* NGSPICE file created from try1.ext - technology: sky130A

X0 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X2 Fvco_By4_QPH_bar.t1 a_66167_26022# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X3 a_28994_17218# a_26368_16652.t2 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X4 a_26690_784.t1 a_23414_5032.t2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X5 Vdd Vso1b a_4226_11420# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X6 a_28220_17218# a_26368_16652.t3 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X7 a_29510_17218# a_26368_16652.t4 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X8 a_23403_5596# a_14188_14050.t2 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X9 a_22629_5596# a_14188_14050.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X10 a_49874_4150.t2 a_49874_4150.t1 a_54950_4814# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.856e+11p ps=1.57e+06u w=1.28e+06u l=8e+06u
X11 a_50320_14126# Fvco_By4_QPH.t2 a_55602_11692# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=1.98421e+11p ps=1.49053e+06u w=1e+06u l=150000u
X12 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X13 vbiasr.t40 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X14 a_29510_17218# a_26368_16652.t5 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X15 a_28994_5597# a_26036_4988.t2 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X16 a_22887_5596# a_14188_14050.t4 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X17 a_54950_4814# a_49874_4150.t4 a_53292_4814# gnd sky130_fd_pr__nfet_01v8 ad=1.856e+11p pd=1.57e+06u as=1.856e+11p ps=1.57e+06u w=1.28e+06u l=8e+06u
X18 a_9354_33563# CLK_BY_4_IPH.t3 vctrl gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=3.012e+11p ps=2.62e+06u w=1e+06u l=150000u
X19 a_26847_11500# a_25099_11445.t2 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X20 Vdd a_66167_26022# a_66154_26414# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X21 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X22 a_24177_5596# a_14188_14050.t5 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X23 gnd a_17685_3840.t17 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X24 a_22629_11500# a_14266_8900.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X25 gnd a_17685_3840.t18 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X26 a_66357_25280# RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=6.405e+10p pd=725000u as=9.2007e+10p ps=682276u w=420000u l=150000u
X27 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X28 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X29 Vdd a_63529_26290# a_63419_26414# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=1.134e+11p ps=1.1e+06u w=420000u l=150000u
X30 a_28736_5597# a_26036_4988.t3 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X31 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X32 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X33 a_26847_11500# a_25099_11445.t3 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X34 a_29510_5597# a_26036_4988.t4 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X35 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X36 gnd Vso3b a_8744_13422# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X37 gnd a_17685_3840.t19 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X38 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X39 gnd Vso5b a_8748_12270# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X40 a_26847_11500# a_25099_11445.t4 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X41 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X42 a_23919_5596# a_14188_14050.t6 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X43 a_28994_5597# a_26036_4988.t5 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X44 a_52052_20860.t9 a_56334_20860.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X45 a_26847_11500# a_25099_11445.t5 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X46 a_23156_5032.t6 a_14188_14050.t7 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X47 a_28736_17218# a_26368_16652.t6 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X48 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X49 a_65546_25646# RESET Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=9.08803e+10p ps=655615u w=420000u l=150000u
X50 a_25299_17217# a_23436_16644.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X51 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X52 a_26847_17217# a_23436_16644.t3 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X53 a_28736_17218# a_26368_16652.t7 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X54 a_25815_5596# a_23414_5032.t3 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X55 a_51276_14152# Fvco_By4_QPH.t3 a_51636_13108# gnd sky130_fd_pr__nfet_01v8 ad=2.07143e+11p pd=1.67714e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X56 gnd a_17685_3840.t20 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X57 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X58 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X59 a_63311_26048# a_62795_26048# a_63216_26048# gnd sky130_fd_pr__nfet_01v8 ad=5.94e+10p pd=690000u as=6.09231e+10p ps=687692u w=360000u l=150000u
X60 vbiasr.t19 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X61 a_23145_5596# a_14188_14050.t8 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X62 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X63 a_26331_11500# a_25099_11445.t6 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X64 a_28478_5597# a_26036_4988.t6 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X65 a_29252_5597# a_26036_4988.t7 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X66 Vdd CLK_IN a_4288_11534# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X67 a_25778_4988.t6 a_23414_5032.t4 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X68 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X69 a_26331_11500# a_25099_11445.t7 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X70 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X71 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X72 gnd a_17685_3840.t21 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X73 a_23145_17217# Fvco.t2 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X74 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X75 a_28220_17218# a_26368_16652.t8 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X76 a_23145_17217# Fvco.t3 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X77 a_52052_20860.t18 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X78 a_56602_11692# vbiasob.t3 a_56272_15934.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=2e+06u
X79 a_27962_5597# a_26036_4988.t8 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X80 vbiasbuffer.t0 a_49874_4150.t5 a_54966_2992# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9575e+11p ps=1.64e+06u w=1.35e+06u l=8e+06u
X81 a_26331_17217# a_23436_16644.t4 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X82 a_28220_17218# a_26368_16652.t9 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X83 vbiasob.t0 a_57726_5786.t5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.23446e+11p ps=1.65695e+06u w=1.02e+06u l=1e+06u
X84 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X85 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X86 a_25557_11500# a_25099_11445.t8 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X87 a_25557_5596# a_23414_5032.t5 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X88 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X89 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X90 gnd gnd vbiasr.t18 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X91 a_22887_5596# a_14188_14050.t9 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X92 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X93 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X94 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X95 a_23661_5596# a_14188_14050.t10 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X96 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X97 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X98 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X99 a_26847_5596# a_23414_5032.t6 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X100 a_28578_5014.t6 a_26036_4988.t9 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X101 gnd gnd vbiasr.t17 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X102 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X103 a_28220_5597# a_26036_4988.t10 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X104 gnd a_17685_3840.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X105 a_24177_11500# a_14266_8900.t3 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X106 a_50583_13108.t0 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X107 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X108 a_25557_11500# a_25099_11445.t9 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X109 a_52052_20860.t8 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X110 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X111 vinit.t39 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X112 a_23403_5596# a_14188_14050.t11 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X113 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X114 a_29252_11501# a_27762_11446.t2 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X115 a_25557_11500# a_25099_11445.t10 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X116 a_25299_5596# a_23414_5032.t7 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X117 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X118 a_49932_4124.t2 a_49932_4124.t1 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=2e+07u
X119 a_28994_5597# a_26036_4988.t11 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X120 a_25557_11500# a_25099_11445.t11 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X121 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X122 a_65438_25280# a_65088_25280# a_65343_25280# Vdd sky130_fd_pr__pfet_01v8_hvt ad=7.245e+10p pd=765000u as=6.51e+10p ps=730000u w=420000u l=150000u
X123 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X124 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X125 a_66346_26048# RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=6.405e+10p pd=725000u as=9.2007e+10p ps=682276u w=420000u l=150000u
X126 a_26589_5596# a_23414_5032.t8 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X127 a_65656_25522# a_65438_25280# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.722e+11p pd=1.58e+06u as=1.81761e+11p ps=1.31123e+06u w=840000u l=150000u
X128 a_24177_11500# a_14266_8900.t4 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X129 vbiasr.t16 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X130 a_44752_16348.t4 a_51138_19904.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X131 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X132 a_25557_17217# a_23436_16644.t5 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X133 vbiasr.t15 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X134 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X135 a_24177_11500# a_14266_8900.t5 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X136 a_27962_11501# a_27762_11446.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X137 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X138 a_14832_12082.t1 a_14188_14050.t12 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X139 a_29252_11501# a_27762_11446.t4 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X140 a_56602_11692# a_51636_13108# a_52052_20860.t17 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X141 a_29510_5597# a_26036_4988.t12 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X142 a_24177_11500# a_14266_8900.t6 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X143 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X144 a_33808_31746# CLK_BY_4_IPH_BAR.t3 a_34044_31208# Vdd sky130_fd_pr__pfet_01v8 ad=3.78914e+11p pd=2.83143e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X145 a_66003_25280# a_64922_25280# a_65656_25522# Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=8.61e+10p ps=790000u w=420000u l=150000u
X146 a_29252_11501# a_27762_11446.t5 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X147 Vdd a_56334_19906# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X148 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X149 a_26073_5596# a_23414_5032.t9 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X150 Vdd Vdd vinit.t38 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X151 a_24177_17217# Fvco.t4 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X152 a_29252_11501# a_27762_11446.t6 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X153 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X154 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X155 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X156 a_26847_17217# a_23436_16644.t6 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X157 a_23160_10936.t6 a_14266_8900.t7 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X158 gnd Vso7b a_8748_11114# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X159 a_29252_17218# a_26368_16652.t10 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X160 a_23661_11500# a_14266_8900.t8 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X161 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X162 a_26847_17217# a_23436_16644.t7 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X163 gnd gnd vbiasr.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X164 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X165 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X166 a_23661_11500# a_14266_8900.t9 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X167 a_25815_5596# a_23414_5032.t10 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X168 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X169 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X170 vinit.t19 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X171 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X172 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X173 a_23919_11500# a_14266_8900.t10 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X174 a_26331_5596# a_23414_5032.t11 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X175 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X176 a_55602_11692# a_51041_13108# a_52052_20860.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X177 a_42574_15624# Fvco_By4_QPH_bar.t2 a_42550_16062# Vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X178 a_29252_5597# a_26036_4988.t13 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X179 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X180 Vdd Vdd vinit.t37 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X181 gnd gnd vbiasr.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X182 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X183 a_53308_3580# a_49874_4150.t6 vbiasr.t20 gnd sky130_fd_pr__nfet_01v8 ad=7.0035e+11p pd=5.12e+06u as=0p ps=0u w=4.83e+06u l=8e+06u
X184 a_23661_17217# Fvco.t5 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X185 a_26331_17217# a_23436_16644.t8 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X186 a_22887_11500# a_14266_8900.t11 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X187 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X188 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X189 CLK_BY_4_IPH_BAR.t1 a_66742_25280# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X190 a_28438_10874.t6 a_27762_11446.t7 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X191 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X192 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X193 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X194 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X195 gnd a_17685_3840.t23 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X196 a_26331_17217# a_23436_16644.t9 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X197 a_23919_11500# a_14266_8900.t12 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X198 gnd a_17685_3840.t24 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X199 a_28438_10874.t5 a_27762_11446.t8 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X200 a_25557_5596# a_23414_5032.t12 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X201 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X202 a_23919_11500# a_14266_8900.t13 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X203 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X204 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X205 a_65438_25280# a_64922_25280# a_65343_25280# gnd sky130_fd_pr__nfet_01v8 ad=5.94e+10p pd=690000u as=6.09231e+10p ps=687692u w=360000u l=150000u
X206 a_23919_11500# a_14266_8900.t14 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X207 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X208 a_63573_26048# a_63529_26290# a_63407_26048# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.50877e+11p ps=1.18462e+06u w=420000u l=150000u
X209 gnd a_17685_3840.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X210 a_22887_11500# a_14266_8900.t15 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X211 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X212 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X213 a_14910_6932.t1 a_14266_8900.t16 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X214 a_28622_16652# a_26368_16652.t11 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X215 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X216 gnd Vso4b a_8740_12844# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X217 a_4314_11564# a_4288_11534# a_4314_11468# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X218 a_23919_17217# Fvco.t4 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X219 a_22887_11500# a_14266_8900.t17 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X220 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X221 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X222 gnd a_17685_3840.t26 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X223 gnd a_17685_3840.t27 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X224 Vdd a_4288_11918# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X225 a_23403_11500# a_14266_8900.t18 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X226 a_22887_11500# a_14266_8900.t19 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X227 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X228 CLK_BY_2_BAR.t0 a_64615_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X229 a_23403_11500# a_14266_8900.t20 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X230 a_26016_10878.t7 a_25099_11445.t12 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X231 a_25299_5596# a_23414_5032.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X232 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X233 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X234 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X235 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X236 a_22887_17217# Fvco.t4 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X237 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X238 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X239 a_64725_25280# CLK_BY_2_BAR.t2 Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.35e+11p pd=1.27e+06u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X240 a_28622_16652# a_26368_16652.t12 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X241 a_25557_17217# a_23436_16644.t10 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X242 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X243 gnd a_17685_3840.t28 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X244 a_25557_17217# a_23436_16644.t11 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X245 a_26073_11500# a_25099_11445.t13 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X246 gnd a_57726_5786.t2 a_57726_5786.t3 gnd sky130_fd_pr__nfet_01v8 ad=6.57193e+11p pd=4.8734e+06u as=0p ps=0u w=3e+06u l=1e+06u
X247 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X248 a_23403_17217# Fvco.t4 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X249 gnd gnd vinit.t18 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X250 a_22629_11500# a_14266_8900.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X251 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X252 a_49932_4124.t0 a_49874_4150.t7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.80402e+11p ps=2.07932e+06u w=1.28e+06u l=8e+06u
X253 a_77280_24640.t1 a_77254_23336.t5 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X254 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X255 a_24177_17217# Fvco.t6 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X256 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X257 a_24177_17217# Fvco.t7 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X258 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X259 gnd RESET a_63573_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=4.41e+10p ps=630000u w=420000u l=150000u
X260 a_29252_17218# a_26368_16652.t13 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X261 vbiasob.t2 vbiasob.t1 a_54448_7822.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X262 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X263 Vso1b a_24410_25128.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X264 a_28478_11501# a_27762_11446.t9 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X265 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X266 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X267 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X268 a_29252_17218# a_26368_16652.t14 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X269 a_22629_11500# a_14266_8900.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X270 a_23308_802.t0 Fvco.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X271 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X272 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X273 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X274 a_26368_16652.t0 a_23436_16644.t12 a_26110_16652# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X275 a_28478_11501# a_27762_11446.t10 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X276 a_24177_5596# a_14188_14050.t13 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X277 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.19064e+11p pd=1.62447e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X278 a_22629_11500# a_14266_8900.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X279 Vdd Vdd vbiasr.t39 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X280 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X281 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X282 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X283 a_22629_11500# a_14266_8900.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X284 a_23661_17217# Fvco.t9 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X285 gnd Vso1b a_8744_9386# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X286 a_28478_17218# a_26368_16652.t15 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X287 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X288 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X289 a_22629_17217# Fvco.t4 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X290 a_23661_17217# Fvco.t10 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X291 a_26036_4988.t0 a_23414_5032.t14 a_17685_3840.t9 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X292 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X293 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X294 Vdd a_4226_11420# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X295 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X296 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X297 gnd a_64725_25280# a_64922_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X298 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X299 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X300 Vdd a_4226_12188# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X301 a_25815_11500# a_25099_11445.t14 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X302 vbiasr.t38 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X303 a_32948_24994.t1 a_27762_11446.t11 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X304 Vso2b a_28790_25040.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X305 vbiasr.t37 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X306 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X307 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X308 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X309 a_28478_17218# a_26368_16652.t16 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X310 a_28622_16652# a_26368_16652.t17 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X311 a_23145_5596# a_14188_14050.t14 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X312 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X313 a_23919_17217# Fvco.t11 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X314 vbiasr.t36 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X315 gnd a_17685_3840.t29 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X316 a_28622_16652# a_26368_16652.t18 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X317 Vdd a_66167_26022# a_66731_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X318 a_23919_17217# Fvco.t12 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X319 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X320 vinit.t17 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X321 a_14910_6932.t0 a_14266_8900.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X322 gnd a_17685_3840.t30 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X323 a_52052_20860.t16 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X324 gnd a_17685_3840.t31 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X325 a_51276_14152# a_51334_14126# a_33808_31746# gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=3.78571e+11p ps=2.99714e+06u w=2e+06u l=1e+06u
X326 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X327 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X328 Vdd a_65992_26048# a_66167_26022# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X329 Vdd Vso6b a_4226_11804# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X330 a_22887_17217# Fvco.t13 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X331 a_29510_11501# a_27762_11446.t12 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X332 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X333 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X334 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X335 a_27962_5597# a_26036_4988.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X336 a_22887_17217# Fvco.t14 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X337 Vdd Vdd vbiasr.t35 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X338 a_51532_4150.t1 a_51532_4150.t0 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.59194e+11p ps=2.59124e+06u w=1.66e+06u l=4e+06u
X339 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X340 Vdd a_65656_25522# a_65546_25646# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=1.134e+11p ps=1.1e+06u w=420000u l=150000u
X341 Vdd CLK_BY_2_BAR.t3 a_64911_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X342 a_56602_11692# a_51636_13108# a_52052_20860.t15 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X343 Vdd a_50032_16080.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X344 a_23403_17217# Fvco.t15 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X345 a_23661_5596# a_14188_14050.t15 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X346 a_22887_5596# a_14188_14050.t16 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X347 a_50511_16072.t7 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X348 Vdd Vdd vinit.t36 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X349 Vdd Vdd vbiasr.t34 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X350 a_64038_26414# a_62961_26048# a_63876_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=5.88e+10p ps=700000u w=420000u l=150000u
X351 a_23403_17217# Fvco.t16 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X352 a_23919_5596# a_14188_14050.t17 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X353 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X354 Vdd a_51138_19904.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X355 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X356 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X357 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X358 a_52052_20860.t6 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X359 a_50583_13108.t1 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X360 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X361 a_65534_25280# a_65088_25280# a_65438_25280# gnd sky130_fd_pr__nfet_01v8 ad=1.29323e+11p pd=1.01538e+06u as=5.94e+10p ps=690000u w=360000u l=150000u
X362 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X363 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X364 a_27962_11501# a_27762_11446.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X365 Vso4b a_38070_8852.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X366 a_52052_20224# a_56272_15934.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X367 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X368 a_14266_8900.t0 a_25099_11445.t15 a_26016_10878.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X369 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X370 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X371 a_28994_5597# a_26036_4988.t15 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X372 Vso5b a_14910_6932.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X373 a_26589_11500# a_25099_11445.t16 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X374 vbiasr.t33 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X375 a_55602_11692# a_51041_13108# a_52052_20860.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X376 a_26589_11500# a_25099_11445.t17 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X377 a_23919_5596# a_14188_14050.t18 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X378 a_24177_5596# a_14188_14050.t19 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X379 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X380 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X381 Fvco_By4_QPH_bar.t0 a_66167_26022# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X382 a_23160_10936.t5 a_14266_8900.t26 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X383 a_27962_11501# a_27762_11446.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X384 a_64230_26048# RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=6.405e+10p pd=725000u as=9.2007e+10p ps=682276u w=420000u l=150000u
X385 a_56602_11692# a_51636_13108# a_52052_20860.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X386 a_27962_11501# a_27762_11446.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X387 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X388 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X389 a_28478_17218# a_26368_16652.t19 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X390 a_30384_802.t1 a_26036_4988.t16 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X391 a_77598_24640.t1 a_77572_23336.t3 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X392 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X393 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X394 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X395 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X396 a_4314_12044# a_4226_11996# a_4314_11948# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X397 a_26589_17217# a_23436_16644.t13 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X398 a_22629_17217# Fvco.t17 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X399 a_27962_11501# a_27762_11446.t16 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X400 gnd CLK_BY_2_BAR.t4 a_64911_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X401 a_65656_25522# a_65438_25280# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.27872e+11p pd=1.2608e+06u as=1.40201e+11p ps=1.03966e+06u w=640000u l=150000u
X402 a_28478_17218# a_26368_16652.t20 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X403 a_26073_5596# a_23414_5032.t15 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X404 a_22629_17217# Fvco.t18 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X405 a_23145_11500# a_14266_8900.t27 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X406 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X407 a_23160_10936.t4 a_14266_8900.t28 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X408 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X409 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X410 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X411 a_27962_17218# a_26368_16652.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X412 a_51041_13108# a_50511_16072.t8 a_50583_13108.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X413 a_66167_26022# RESET Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X414 a_23160_10936.t3 a_14266_8900.t29 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X415 a_28220_11501# a_27762_11446.t17 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X416 a_28578_5014.t5 a_26036_4988.t17 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X417 a_57726_5786.t4 a_51532_4150.t4 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.72176e+11p ps=2.6849e+06u w=1.72e+06u l=4e+06u
X418 a_23160_10936.t2 a_14266_8900.t30 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X419 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X420 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X421 a_26847_17217# a_23436_16644.t14 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X422 a_63311_26048# a_62961_26048# a_63216_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=7.245e+10p pd=765000u as=6.51e+10p ps=730000u w=420000u l=150000u
X423 a_55602_11692# a_51041_13108# a_52052_20860.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X424 vinit.t35 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X425 a_65088_25280# a_64922_25280# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X426 a_23403_5596# a_14188_14050.t20 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X427 Vdd a_54410_8156# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X428 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X429 a_23178_16644# Fvco.t19 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X430 CLK_IN a_23308_802.t2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X431 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X432 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X433 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X434 a_50128_8156# a_54448_7822.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X435 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X436 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X437 a_65546_25646# a_64922_25280# a_65438_25280# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=7.245e+10p ps=765000u w=420000u l=150000u
X438 gnd a_17685_3840.t32 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X439 a_53308_2992# a_49874_4150.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.9575e+11p pd=1.64e+06u as=2.95737e+11p ps=2.19303e+06u w=1.35e+06u l=8e+06u
X440 gnd a_17685_3840.t33 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X441 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X442 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X443 a_28578_5014.t4 a_26036_4988.t18 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X444 gnd Vso2b a_8736_14034# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X445 a_27962_5597# a_26036_4988.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X446 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X447 Vdd a_4226_11996# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X448 vbiasr.t12 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X449 gnd a_17685_3840.t34 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X450 Fvco.t0 a_26036_4988.t20 a_28578_5014.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X451 a_22629_5596# a_14188_14050.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X452 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X453 a_26016_10878.t6 a_25099_11445.t18 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X454 a_25299_11500# a_25099_11445.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X455 a_29510_5597# a_26036_4988.t21 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X456 a_23403_5596# a_14188_14050.t22 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X457 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X458 a_17685_3840.t8 vinit.t40 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=1e+06u
X459 a_23661_5596# a_14188_14050.t23 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X460 Vdd a_63876_26048# a_64051_26022# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X461 a_25299_11500# a_25099_11445.t20 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X462 a_23919_5596# a_14188_14050.t24 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X463 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X464 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X465 gnd a_17685_3840.t35 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X466 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X467 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X468 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X469 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X470 a_26073_11500# a_25099_11445.t21 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X471 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X472 a_65077_26048# a_64911_26048# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.38484e+11p ps=999033u w=640000u l=150000u
X473 a_25299_17217# a_23436_16644.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X474 Vso7b a_26690_784.t2 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X475 a_30384_802.t0 a_26036_4988.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X476 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X477 a_26016_10878.t5 a_25099_11445.t22 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X478 a_25815_5596# a_23414_5032.t16 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X479 a_28736_5597# a_26036_4988.t23 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X480 a_26016_10878.t4 a_25099_11445.t23 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X481 a_29252_5597# a_26036_4988.t24 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X482 a_29510_5597# a_26036_4988.t25 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X483 a_66112_25280# a_64922_25280# a_66003_25280# gnd sky130_fd_pr__nfet_01v8 ad=6.17538e+10p pd=692308u as=7.11e+10p ps=755000u w=360000u l=150000u
X484 a_26016_10878.t3 a_25099_11445.t24 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X485 gnd a_17685_3840.t36 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X486 a_26073_11500# a_25099_11445.t25 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X487 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X488 a_56602_11692# Fvco_By4_QPH_bar.t3 a_50320_14126# gnd sky130_fd_pr__nfet_01v8 ad=1.98421e+11p pd=1.49053e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X489 a_23156_5032.t5 a_14188_14050.t25 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X490 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X491 gnd a_17685_3840.t37 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X492 a_46856_21176.t1 a_51138_21494.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X493 gnd a_17685_3840.t38 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X494 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X495 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X496 a_26110_16652# a_23436_16644.t16 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X497 a_25557_17217# a_23436_16644.t17 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X498 a_26073_11500# a_25099_11445.t26 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X499 a_65645_26290# a_65427_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.27872e+11p pd=1.2608e+06u as=1.40201e+11p ps=1.03966e+06u w=640000u l=150000u
X500 a_26589_17217# a_23436_16644.t18 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X501 a_77280_24640.t2 a_77254_23336.t4 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X502 a_26073_11500# a_25099_11445.t27 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X503 vbiasr.t11 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X504 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X505 a_26589_17217# a_23436_16644.t19 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X506 a_25815_5596# a_23414_5032.t17 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X507 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X508 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X509 a_27962_17218# a_26368_16652.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X510 a_25557_5596# a_23414_5032.t18 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X511 a_42574_15624# vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=4e+06u
X512 gnd a_56334_20860.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X513 a_26073_5596# a_23414_5032.t19 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X514 a_28478_5597# a_26036_4988.t26 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X515 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X516 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X517 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X518 gnd a_64051_26022# a_64615_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X519 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X520 a_29252_5597# a_26036_4988.t27 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X521 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X522 a_26073_17217# a_23436_16644.t20 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X523 a_24177_17217# Fvco.t20 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X524 a_27962_17218# a_26368_16652.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X525 a_25778_4988.t5 a_23414_5032.t20 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X526 gnd a_17685_3840.t39 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X527 a_26331_11500# a_25099_11445.t28 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X528 gnd gnd vinit.t16 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X529 Vdd vinit.t41 a_17685_3840.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=2.16382e+11p pd=1.56099e+06u as=0p ps=0u w=1e+06u l=1e+06u
X530 a_28578_5014.t3 a_26036_4988.t28 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X531 a_65077_26048# a_64911_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X532 Vdd Vso3b a_4288_12110# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X533 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X534 Vdd CLK_BY_2_BAR.t5 a_64725_25280# Vdd sky130_fd_pr__pfet_01v8_hvt ad=2.16382e+11p pd=1.56099e+06u as=1.35e+11p ps=1.27e+06u w=1e+06u l=150000u
X535 Vdd Vso5b a_4288_11918# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X536 a_23178_16644# Fvco.t21 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X537 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X538 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X539 a_34044_31208# CLK_BY_4_IPH.t4 a_33808_31746# gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=1.89286e+11p ps=1.49857e+06u w=1e+06u l=150000u
X540 Vso3b a_32948_24994.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X541 a_25815_11500# a_25099_11445.t29 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X542 gnd gnd vbiasr.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X543 a_23403_5596# a_14188_14050.t26 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X544 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X545 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X546 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X547 a_23178_16644# Fvco.t22 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X548 a_25557_5596# a_23414_5032.t21 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X549 a_23504_23306# Vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X550 a_25299_5596# a_23414_5032.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X551 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X552 a_33808_31746# CLK_BY_4_IPH_BAR.t4 a_9354_33563# gnd sky130_fd_pr__nfet_01v8 ad=1.89286e+11p pd=1.49857e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X553 a_51636_13108# a_50511_16072.t9 a_46856_19268.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X554 a_77280_24640.t0 CLK_BY_4_IPH_BAR.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X555 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X556 a_26847_5596# a_23414_5032.t23 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X557 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X558 a_25815_11500# a_25099_11445.t30 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X559 bb Fvco_By4_QPH.t4 a_47968_16078# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X560 a_28220_5597# a_26036_4988.t29 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X561 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X562 Vdd Vdd vinit.t34 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X563 Vdd Vso7b a_4226_11612# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X564 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X565 a_29510_11501# a_27762_11446.t18 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X566 a_25815_11500# a_25099_11445.t31 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X567 a_29510_5597# a_26036_4988.t30 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X568 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X569 a_25815_11500# a_25099_11445.t32 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X570 a_47968_16078# Fvco_By4_QPH_bar.t4 aa Vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X571 a_25299_5596# a_23414_5032.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X572 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X573 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X574 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X575 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X576 Vso3b a_32948_24994.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X577 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X578 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X579 Vdd Vso7b a_4288_11726# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X580 a_25815_17217# a_23436_16644.t21 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X581 a_25299_17217# a_23436_16644.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X582 a_26589_5596# a_23414_5032.t25 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X583 a_23919_17217# Fvco.t23 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X584 a_9354_33563# CLK_BY_4_IPH.t5 a_33808_31746# Vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.78914e+11p ps=2.83143e+06u w=2e+06u l=150000u
X585 a_25299_17217# a_23436_16644.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X586 a_29510_11501# a_27762_11446.t19 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X587 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X588 a_25815_5596# a_23414_5032.t26 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X589 a_63407_26048# a_62961_26048# a_63311_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.29323e+11p pd=1.01538e+06u as=5.94e+10p ps=690000u w=360000u l=150000u
X590 a_29510_11501# a_27762_11446.t20 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X591 CLK_IN a_23308_802.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X592 a_66101_26048# a_64911_26048# a_65992_26048# gnd sky130_fd_pr__nfet_01v8 ad=6.17538e+10p pd=692308u as=7.11e+10p ps=755000u w=360000u l=150000u
X593 a_25099_11445.t0 a_27762_11446.t21 a_28438_10874.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X594 a_28790_25040.t1 a_26368_16652.t24 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X595 a_22887_17217# Fvco.t24 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X596 a_29510_11501# a_27762_11446.t22 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X597 a_29252_5597# a_26036_4988.t31 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X598 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X599 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X600 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X601 a_65535_26414# RESET Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=9.08803e+10p ps=655615u w=420000u l=150000u
X602 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X603 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X604 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X605 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X606 a_26110_16652# a_23436_16644.t24 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X607 Vso5b a_14910_6932.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X608 a_23436_16644.t0 Fvco.t4 a_17685_3840.t5 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X609 vbiasot vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=4e+06u
X610 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X611 a_29510_17218# a_26368_16652.t25 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X612 Vso7b a_26690_784.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X613 a_26110_16652# a_23436_16644.t25 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X614 a_77598_24640.t2 a_77572_23336.t2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X615 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X616 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X617 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X618 a_23661_11500# a_14266_8900.t31 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X619 a_26073_17217# a_23436_16644.t26 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X620 a_25557_5596# a_23414_5032.t27 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X621 Vdd Vso8b a_4288_11534# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X622 a_26331_5596# a_23414_5032.t28 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X623 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X624 gnd a_17685_3840.t40 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X625 a_26073_17217# a_23436_16644.t27 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X626 gnd a_17685_3840.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X627 a_50262_14152# Fvco_By4_QPH.t5 a_51041_13108# gnd sky130_fd_pr__nfet_01v8 ad=2.07143e+11p pd=1.67714e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X628 a_47968_16078# a_42550_16062# a_50511_16072.t1 Vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X629 CLK_BY_2 a_64051_26022# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X630 a_23145_11500# a_14266_8900.t32 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X631 a_49874_4150.t0 a_51532_4150.t5 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.59194e+11p ps=2.59124e+06u w=1.66e+06u l=4e+06u
X632 Vdd CLK_IN a_4226_11420# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X633 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X634 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X635 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X636 bb vbiasbuffer.t3 a_51826_16054.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=1e+06u
X637 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X638 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X639 a_28220_11501# a_27762_11446.t23 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X640 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X641 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X642 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.0669e+12p pd=2.27425e+07u as=3.0669e+12p ps=2.27425e+07u w=1.4e+07u l=1e+06u
X643 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X644 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X645 a_28438_10874.t4 a_27762_11446.t24 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X646 a_43010_16058# Fvco_By4_QPH.t6 a_42574_15624# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X647 a_25299_5596# a_23414_5032.t29 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X648 Fvco_By4_QPH.t1 a_66731_26048# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X649 a_28994_11501# a_27762_11446.t25 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X650 a_23145_11500# a_14266_8900.t33 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X651 Vdd Vdd vbiasr.t32 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X652 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X653 a_22629_17217# Fvco.t25 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X654 a_28994_11501# a_27762_11446.t26 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X655 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X656 a_23145_11500# a_14266_8900.t34 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X657 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X658 a_28220_11501# a_27762_11446.t27 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X659 a_23145_11500# a_14266_8900.t35 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X660 a_50511_16072.t6 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X661 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X662 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X663 a_66165_25646# a_65088_25280# a_66003_25280# Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=5.88e+10p ps=700000u w=420000u l=150000u
X664 a_28220_11501# a_27762_11446.t28 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X665 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X666 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X667 a_64051_26022# RESET Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X668 a_65427_26048# a_65077_26048# a_65332_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=7.245e+10p pd=765000u as=6.51e+10p ps=730000u w=420000u l=150000u
X669 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X670 Vdd Vdd vinit.t33 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X671 a_17685_3840.t1 vinit.t42 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=1e+06u
X672 a_23145_17217# Fvco.t4 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X673 a_28994_17218# a_26368_16652.t26 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X674 a_28220_11501# a_27762_11446.t29 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X675 a_42782_16060# vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=4e+06u
X676 Vdd a_51138_19904.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X677 a_77598_24640.t0 CLK_BY_4_IPH.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X678 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X679 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X680 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X681 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X682 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X683 a_25815_17217# a_23436_16644.t28 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X684 a_23403_11500# a_14266_8900.t36 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X685 a_28220_17218# a_26368_16652.t27 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X686 a_25815_17217# a_23436_16644.t29 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X687 vinit.t15 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X688 vctrl CLK_BY_4_IPH_BAR.t5 a_34044_31208# gnd sky130_fd_pr__nfet_01v8 ad=3.012e+11p pd=2.62e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X689 a_65992_26048# a_64911_26048# a_65645_26290# Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=8.61e+10p ps=790000u w=420000u l=150000u
X690 a_52052_20224# a_56334_19906# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X691 a_28994_17218# a_26368_16652.t28 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X692 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X693 a_24177_5596# a_14188_14050.t27 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X694 a_42550_16062# Fvco_By4_QPH.t7 a_42574_15624# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X695 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X696 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X697 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X698 a_23436_16644.t1 Fvco.t26 a_23178_16644# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X699 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X700 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X701 a_29510_17218# a_26368_16652.t29 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X702 a_22629_5596# a_14188_14050.t28 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X703 Vdd Vdd vbiasr.t31 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X704 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X705 a_66003_25280# a_65088_25280# a_65656_25522# gnd sky130_fd_pr__nfet_01v8 ad=7.11e+10p pd=755000u as=7.1928e+10p ps=709200u w=360000u l=150000u
X706 Vso6b a_14832_12082.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X707 a_28736_11501# a_27762_11446.t30 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X708 gnd a_17685_3840.t42 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X709 a_4314_11660# a_4226_11612# a_4314_11564# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X710 a_29510_17218# a_26368_16652.t30 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X711 gnd a_17685_3840.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X712 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X713 a_65343_25280# CLK_BY_4_IPH_BAR.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=7.10769e+10p pd=802308u as=9.2007e+10p ps=682276u w=420000u l=150000u
X714 a_28736_11501# a_27762_11446.t31 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X715 a_23919_5596# a_14188_14050.t29 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X716 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X717 a_28478_11501# a_27762_11446.t32 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X718 a_24177_5596# a_14188_14050.t30 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X719 a_23414_5032.t1 a_14188_14050.t31 a_17685_3840.t11 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X720 Vdd Vdd vinit.t32 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X721 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X722 vinit.t31 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X723 Vdd vinit.t43 a_17685_3840.t2 Vdd sky130_fd_pr__pfet_01v8_lvt ad=2.16382e+11p pd=1.56099e+06u as=0p ps=0u w=1e+06u l=1e+06u
X724 a_28736_17218# a_26368_16652.t31 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X725 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X726 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X727 gnd a_17685_3840.t44 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X728 a_28736_5597# a_26036_4988.t32 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X729 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X730 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X731 gnd a_17685_3840.t45 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X732 gnd a_17685_3840.t46 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X733 a_26331_11500# a_25099_11445.t33 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X734 a_23156_5032.t4 a_14188_14050.t32 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X735 a_77572_23336.t5 a_77254_23336.t1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X736 Vdd Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X737 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X738 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X739 vbiasr.t30 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X740 vbiasr.t29 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X741 a_28736_17218# a_26368_16652.t32 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X742 a_27962_5597# a_26036_4988.t33 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X743 vinit.t14 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X744 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X745 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X746 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X747 a_4314_11756# a_4288_11726# a_4314_11660# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X748 a_28478_5597# a_26036_4988.t34 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X749 a_23145_5596# a_14188_14050.t33 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X750 gnd gnd vinit.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X751 a_26331_11500# a_25099_11445.t34 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X752 a_23661_5596# a_14188_14050.t34 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X753 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X754 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X755 a_25778_4988.t4 a_23414_5032.t30 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X756 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X757 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X758 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X759 a_28994_17218# a_26368_16652.t33 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X760 a_26331_11500# a_25099_11445.t35 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X761 a_28578_5014.t2 a_26036_4988.t35 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X762 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X763 a_23145_17217# Fvco.t27 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X764 a_23308_802.t1 Fvco.t28 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X765 a_28994_17218# a_26368_16652.t34 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X766 a_26331_11500# a_25099_11445.t36 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X767 a_23145_17217# Fvco.t29 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X768 a_42782_16060# Fvco_By4_QPH_bar.t5 a_43010_16058# Vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X769 a_27962_5597# a_26036_4988.t36 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X770 a_28220_17218# a_26368_16652.t35 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X771 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X772 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X773 a_65343_25280# CLK_BY_4_IPH_BAR.t7 Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=6.51e+10p pd=730000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X774 CLK_BY_4_IPH.t1 a_66178_25254# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X775 a_26331_17217# a_23436_16644.t30 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X776 a_23403_5596# a_14188_14050.t35 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X777 vinit.t30 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X778 a_23178_16644# Fvco.t30 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X779 a_28220_17218# a_26368_16652.t36 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X780 Vdd Vdd vbiasr.t28 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X781 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X782 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X783 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X784 a_22887_5596# a_14188_14050.t36 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X785 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X786 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X787 gnd a_17685_3840.t47 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X788 a_23661_5596# a_14188_14050.t37 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X789 a_26847_5596# a_23414_5032.t31 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X790 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X791 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X792 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X793 Vdd Vso8b a_4226_11612# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X794 vbiasr.t9 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X795 a_24177_5596# a_14188_14050.t38 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X796 vinit.t29 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X797 a_65992_26048# a_65077_26048# a_65645_26290# gnd sky130_fd_pr__nfet_01v8 ad=7.11e+10p pd=755000u as=7.1928e+10p ps=709200u w=360000u l=150000u
X798 a_28220_5597# a_26036_4988.t37 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X799 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X800 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X801 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X802 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X803 Vdd Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X804 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X805 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X806 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X807 a_65332_26048# Fvco_By4_QPH.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=7.10769e+10p pd=802308u as=9.2007e+10p ps=682276u w=420000u l=150000u
X808 vbiasr.t8 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X809 a_46856_19268.t0 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X810 a_23414_5032.t0 a_14188_14050.t39 a_23156_5032.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X811 a_22629_5596# a_14188_14050.t40 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X812 a_26847_11500# a_25099_11445.t37 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X813 a_29510_5597# a_26036_4988.t38 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X814 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X815 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X816 Vdd Vso6b a_4288_11726# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X817 a_26073_5596# a_23414_5032.t32 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X818 a_46856_21176.t0 a_51138_20858# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X819 a_26847_11500# a_25099_11445.t38 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X820 a_28994_5597# a_26036_4988.t39 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X821 a_26589_11500# a_25099_11445.t39 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X822 a_51826_16054.t1 Vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X823 a_26589_5596# a_23414_5032.t33 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X824 a_26036_4988.t1 a_23414_5032.t14 a_25778_4988.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X825 gnd gnd vinit.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X826 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X827 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X828 a_28736_17218# a_26368_16652.t37 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X829 gnd gnd vbiasr.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X830 gnd a_56334_20860.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X831 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X832 a_26847_17217# a_23436_16644.t31 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X833 a_28736_17218# a_26368_16652.t38 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X834 a_14266_8900.t1 a_25099_11445.t40 a_17685_3840.t6 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X835 a_23661_11500# a_14266_8900.t37 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X836 a_25815_5596# a_23414_5032.t34 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X837 a_51636_13108# Fvco_By4_QPH_bar.t6 a_51276_14152# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X838 a_28736_5597# a_26036_4988.t40 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X839 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X840 a_29252_5597# a_26036_4988.t41 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X841 gnd gnd vbiasr.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X842 gnd gnd vbiasr.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X843 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X844 bb Fvco_By4_QPH.t9 a_47760_15642# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X845 a_26073_5596# a_23414_5032.t35 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X846 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X847 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X848 a_38070_8852.t0 a_25099_11445.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X849 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X850 Vdd Vso2b a_4226_12188# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X851 a_23156_5032.t3 a_14188_14050.t41 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X852 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X853 a_26110_16652# a_23436_16644.t32 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X854 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X855 a_23661_11500# a_14266_8900.t38 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X856 a_27962_5597# a_26036_4988.t42 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X857 Vdd Vdd vinit.t28 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X858 a_23661_11500# a_14266_8900.t39 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X859 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X860 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X861 a_28438_10874.t3 a_27762_11446.t33 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X862 a_26331_5596# a_23414_5032.t36 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X863 a_25557_5596# a_23414_5032.t37 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X864 a_55602_11692# Fvco_By4_QPH_bar.t7 a_50320_14126# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X865 gnd a_17685_3840.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X866 a_28478_5597# a_26036_4988.t43 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X867 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X868 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X869 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X870 a_23661_11500# a_14266_8900.t40 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X871 vbiasr.t4 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X872 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X873 a_23661_5596# a_14188_14050.t42 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X874 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X875 Vdd Vso3b a_4226_11996# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X876 a_26073_17217# a_23436_16644.t33 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X877 a_27762_11446.t1 a_26368_16652.t39 a_28622_16652# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X878 gnd a_17685_3840.t49 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X879 a_25778_4988.t3 a_23414_5032.t38 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X880 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X881 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X882 a_57726_5786.t1 a_57726_5786.t0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.57193e+11p ps=4.8734e+06u w=3e+06u l=1e+06u
X883 Vdd Vdd vinit.t27 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X884 Vdd a_65645_26290# a_65535_26414# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=1.134e+11p ps=1.1e+06u w=420000u l=150000u
X885 a_8752_10532# Vso7b a_4226_11612# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X886 a_23661_17217# Fvco.t4 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X887 aa Fvco_By4_QPH.t10 a_47968_16078# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X888 a_4314_12140# a_4288_12110# a_4314_12044# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X889 a_26331_17217# a_23436_16644.t34 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X890 a_28438_10874.t2 a_27762_11446.t34 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X891 a_56602_11692# a_51636_13108# a_52052_20860.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X892 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X893 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X894 a_25557_11500# a_25099_11445.t42 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X895 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X896 a_62961_26048# a_62795_26048# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.38484e+11p ps=999033u w=640000u l=150000u
X897 gnd a_17685_3840.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X898 a_26331_17217# a_23436_16644.t35 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X899 a_28438_10874.t1 a_27762_11446.t35 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X900 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X901 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X902 gnd gnd vinit.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X903 a_25557_11500# a_25099_11445.t43 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X904 Fvco.t1 a_26036_4988.t44 a_17685_3840.t15 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X905 a_25299_5596# a_23414_5032.t39 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X906 a_23403_11500# a_14266_8900.t41 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X907 a_28438_10874.t0 a_27762_11446.t36 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X908 a_55602_11692# Fvco_By4_QPH_bar.t8 a_51334_14126# gnd sky130_fd_pr__nfet_01v8 ad=1.98421e+11p pd=1.49053e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X909 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X910 a_25299_11500# a_25099_11445.t44 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X911 gnd gnd vbiasr.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X912 Vdd a_66178_25254# a_66742_25280# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X913 a_26847_5596# a_23414_5032.t40 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X914 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X915 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X916 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X917 a_28622_16652# a_26368_16652.t40 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X918 a_25557_17217# a_23436_16644.t36 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X919 a_24177_11500# a_14266_8900.t42 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X920 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X921 a_28220_5597# a_26036_4988.t45 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X922 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X923 a_26690_784.t0 a_23414_5032.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X924 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X925 a_29252_11501# a_27762_11446.t37 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X926 a_24177_11500# a_14266_8900.t43 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X927 a_23403_11500# a_14266_8900.t44 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X928 a_77598_24640.t3 a_77572_23336.t1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X929 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X930 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X931 a_29252_11501# a_27762_11446.t38 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X932 a_55602_11692# a_51041_13108# a_52052_20860.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X933 a_26073_5596# a_23414_5032.t42 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X934 a_23403_11500# a_14266_8900.t45 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X935 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X936 a_54966_3580# a_49874_4150.t9 a_53308_3580# gnd sky130_fd_pr__nfet_01v8 ad=7.0035e+11p pd=5.12e+06u as=7.0035e+11p ps=5.12e+06u w=4.83e+06u l=8e+06u
X937 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X938 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X939 a_24177_17217# Fvco.t31 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X940 a_23403_11500# a_14266_8900.t46 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X941 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X942 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X943 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X944 a_25815_17217# a_23436_16644.t37 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X945 a_47760_15642# Fvco_By4_QPH_bar.t9 bb Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.33143e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X946 a_26589_5596# a_23414_5032.t43 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X947 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X948 a_63216_26048# CLK_BY_2_BAR.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=7.10769e+10p pd=802308u as=9.2007e+10p ps=682276u w=420000u l=150000u
X949 a_26847_17217# a_23436_16644.t38 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X950 a_14188_14050.t1 a_14266_8900.t47 a_23160_10936.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X951 vinit.t26 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X952 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X953 gnd a_4226_12188# a_4314_12140# gnd sky130_fd_pr__nfet_01v8 ad=7.09769e+11p pd=5.26327e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X954 Vdd Vso5b a_4226_11804# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X955 a_29252_17218# a_26368_16652.t41 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X956 a_23403_17217# Fvco.t4 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X957 a_26847_17217# a_23436_16644.t39 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X958 a_28478_11501# a_27762_11446.t39 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X959 a_51334_14126# Fvco_By4_QPH.t11 a_55602_11692# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X960 a_62961_26048# a_62795_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X961 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X962 Vdd a_64051_26022# a_64615_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X963 gnd a_17685_3840.t51 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X964 Vdd a_66178_25254# a_66165_25646# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X965 vinit.t25 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X966 vinit.t10 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X967 Vso2b a_28790_25040.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X968 a_65700_25280# a_65656_25522# a_65534_25280# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.50877e+11p ps=1.18462e+06u w=420000u l=150000u
X969 a_29252_17218# a_26368_16652.t42 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X970 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X971 a_47760_15642# Fvco_By4_QPH_bar.t10 aa gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X972 a_22972_23306.t0 a_23504_23306# gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X973 a_28478_11501# a_27762_11446.t40 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X974 a_50262_14152# a_50320_14126# a_50511_16072.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X975 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X976 Vdd CLK_IN a_62795_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X977 CLK_BY_4_IPH_BAR.t0 a_66742_25280# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X978 a_23919_11500# a_14266_8900.t48 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X979 a_28478_11501# a_27762_11446.t41 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X980 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X981 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X982 a_65535_26414# a_64911_26048# a_65427_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=7.245e+10p ps=765000u w=420000u l=150000u
X983 Vdd a_54468_7504.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X984 a_23919_11500# a_14266_8900.t49 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X985 a_28478_11501# a_27762_11446.t42 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X986 a_26331_5596# a_23414_5032.t44 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X987 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X988 a_23661_17217# Fvco.t32 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X989 a_22887_11500# a_14266_8900.t50 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X990 a_47968_16078# Fvco_By4_QPH_bar.t11 bb gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X991 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X992 Vso1b a_24410_25128.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X993 a_28478_17218# a_26368_16652.t43 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X994 a_23661_17217# Fvco.t33 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X995 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X996 a_23919_17217# Fvco.t34 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X997 a_22887_11500# a_14266_8900.t51 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X998 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X999 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1000 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1001 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1002 vinit.t24 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1003 a_42550_16062# Fvco_By4_QPH.t12 a_42782_16060# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X1004 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1005 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1006 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1007 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1008 a_22887_17217# Fvco.t4 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1009 Vso4b a_38070_8852.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1010 a_52052_20860.t12 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X1011 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1012 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1013 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1014 CLK_BY_2 a_64051_26022# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X1015 a_28622_16652# a_26368_16652.t44 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1016 a_23145_5596# a_14188_14050.t43 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1017 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1018 gnd RESET a_65700_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=4.41e+10p ps=630000u w=420000u l=150000u
X1019 gnd a_66178_25254# a_66112_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=7.20462e+10p ps=807692u w=420000u l=150000u
X1020 a_25557_17217# a_23436_16644.t40 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1021 a_51532_4150.t3 a_49932_4124.t3 a_49874_4150.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.28e+06u l=8e+06u
X1022 Vdd Vdd vbiasr.t27 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1023 Vdd Vdd vbiasr.t26 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1024 a_64725_25280# CLK_BY_2_BAR.t7 gnd gnd sky130_fd_pr__nfet_01v8 ad=8.775e+10p pd=920000u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X1025 Vdd a_4288_11534# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1026 a_28622_16652# a_26368_16652.t45 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1027 CLK_BY_4_IPH.t2 a_66178_25254# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X1028 a_17685_3840.t14 vctrl a_22972_23306.t4 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1029 a_25557_17217# a_23436_16644.t41 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1030 gnd CLK_IN a_62795_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1031 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1032 a_77280_24640.t3 a_77254_23336.t3 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1033 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1034 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1035 a_23145_17217# Fvco.t35 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1036 a_24177_17217# Fvco.t36 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1037 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1038 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1039 gnd a_17685_3840.t52 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1040 Vdd Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1041 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1042 a_24177_17217# Fvco.t37 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1043 gnd a_17685_3840.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1044 a_29252_17218# a_26368_16652.t46 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1045 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1046 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1047 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1048 a_65645_26290# a_65427_26048# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.722e+11p pd=1.58e+06u as=1.81761e+11p ps=1.31123e+06u w=840000u l=150000u
X1049 a_23403_17217# Fvco.t38 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1050 a_22887_5596# a_14188_14050.t44 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1051 vbiasr.t25 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1052 a_52052_20860.t2 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X1053 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1054 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1055 a_29252_17218# a_26368_16652.t47 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1056 a_23403_17217# Fvco.t39 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1057 a_26589_11500# a_25099_11445.t45 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1058 a_22629_11500# a_14266_8900.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1059 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1060 a_24177_5596# a_14188_14050.t45 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1061 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1062 a_22629_11500# a_14266_8900.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1063 vbiasr.t24 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1064 a_50511_16072.t0 a_42550_16062# a_47968_16078# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1065 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1066 Vdd a_51138_20858# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1067 gnd a_17685_3840.t54 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1068 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1069 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1070 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1071 a_22629_17217# Fvco.t4 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1072 vinit.t9 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1073 Fvco_By4_QPH.t0 a_66731_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X1074 Vso6b a_14832_12082.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1075 Vdd Vso4b a_4226_11996# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1076 a_26589_11500# a_25099_11445.t46 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1077 a_28994_5597# a_26036_4988.t46 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1078 a_56602_11692# a_51636_13108# a_52052_20860.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1079 a_50511_16072.t4 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1080 a_51276_14152# Fvco_By4_QPH.t13 a_51041_13108# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1081 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1082 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1083 a_26589_11500# a_25099_11445.t47 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1084 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1085 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1086 a_26589_11500# a_25099_11445.t48 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1087 Vdd Vdd vbiasr.t23 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1088 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1089 a_28478_17218# a_26368_16652.t48 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1090 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1091 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1092 a_34044_31208# CLK_BY_4_IPH.t6 vctrl Vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X1093 Vdd Vso1b a_4226_12188# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1094 a_26589_17217# a_23436_16644.t42 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1095 a_23919_17217# Fvco.t40 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1096 a_28478_17218# a_26368_16652.t49 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1097 a_28994_11501# a_27762_11446.t43 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1098 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1099 a_56602_11692# Fvco_By4_QPH_bar.t12 a_51334_14126# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1100 a_63419_26414# a_62795_26048# a_63311_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=7.245e+10p ps=765000u w=420000u l=150000u
X1101 a_23919_17217# Fvco.t41 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1102 a_43010_16058# Fvco_By4_QPH.t14 a_42782_16060# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1103 a_55602_11692# a_51041_13108# a_52052_20860.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1104 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1105 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1106 vctrl CLK_BY_4_IPH_BAR.t8 a_9354_33563# Vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X1107 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1108 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1109 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1110 a_24410_25128.t0 a_23436_16644.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1111 a_63876_26048# a_62795_26048# a_63529_26290# Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=8.61e+10p ps=790000u w=420000u l=150000u
X1112 a_22887_17217# Fvco.t42 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1113 a_27962_5597# a_26036_4988.t47 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1114 a_53292_4814# a_49874_4150.t10 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.856e+11p pd=1.57e+06u as=2.80402e+11p ps=2.07932e+06u w=1.28e+06u l=8e+06u
X1115 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1116 gnd a_66167_26022# a_66101_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=7.20462e+10p ps=807692u w=420000u l=150000u
X1117 gnd RESET a_65689_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=4.41e+10p ps=630000u w=420000u l=150000u
X1118 a_22887_17217# Fvco.t43 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1119 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1120 vbiasr.t22 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1121 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1122 gnd a_17685_3840.t55 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1123 a_22629_5596# a_14188_14050.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1124 gnd a_17685_3840.t56 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1125 a_23145_5596# a_14188_14050.t47 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1126 a_63529_26290# a_63311_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.27872e+11p pd=1.2608e+06u as=1.40201e+11p ps=1.03966e+06u w=640000u l=150000u
X1127 a_23661_5596# a_14188_14050.t48 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1128 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.0669e+12p pd=2.27425e+07u as=3.0669e+12p ps=2.27425e+07u w=1.4e+07u l=1e+06u
X1129 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.19064e+11p pd=1.62447e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1130 b.t0 a_77572_23336.t4 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1131 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1132 a_28790_25040.t0 a_26368_16652.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1133 a_25299_11500# a_25099_11445.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1134 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1135 vinit.t8 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1136 Vso8b a_30384_802.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X1137 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1138 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1139 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1140 Vdd Vso2b a_4288_12110# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1141 a_46856_19268.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1142 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1143 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1144 Vdd Vso4b a_4288_11918# Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1145 a_56602_11692# a_51636_13108# a_52052_20860.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1146 gnd a_17685_3840.t57 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1147 a_42782_16060# bb a_44752_16348.t3 Vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1148 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1149 a_64051_26022# a_63876_26048# a_64230_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=6.405e+10p ps=725000u w=420000u l=150000u
X1150 a_8748_11114# Vso6b a_4288_11726# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1151 a_26331_17217# a_23436_16644.t44 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1152 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1153 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1154 a_28736_5597# a_26036_4988.t48 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1155 a_22629_5596# a_14188_14050.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1156 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1157 a_25299_11500# a_25099_11445.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1158 a_22887_5596# a_14188_14050.t50 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1159 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1160 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1161 a_25299_11500# a_25099_11445.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1162 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1163 a_23919_5596# a_14188_14050.t51 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1164 a_28736_11501# a_27762_11446.t44 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1165 vbiasot a_51532_4150.t6 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.566e+11p pd=1.66e+06u as=1.16846e+11p ps=842934u w=540000u l=8e+06u
X1166 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1167 a_27962_11501# a_27762_11446.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1168 a_25299_11500# a_25099_11445.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1169 a_23156_5032.t2 a_14188_14050.t52 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1170 vbiasbuffer.t2 vbiasbuffer.t1 a_54468_7504.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1171 a_77572_23336.t6 a_77254_23336.t0 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1172 a_14188_14050.t0 a_14266_8900.t54 a_17685_3840.t4 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1173 a_27962_11501# a_27762_11446.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1174 a_55602_11692# a_51041_13108# a_52052_20860.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1175 a_51334_14126# Fvco_By4_QPH.t15 a_56602_11692# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=1.98421e+11p ps=1.49053e+06u w=1e+06u l=150000u
X1176 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1177 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1178 a_25299_17217# a_23436_16644.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1179 a_22629_17217# Fvco.t44 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1180 vbiasr.t2 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1181 gnd a_17685_3840.t58 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1182 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1183 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1184 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1185 a_42574_15624# aa a_44752_16348.t1 Vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1186 a_26073_5596# a_23414_5032.t45 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1187 a_28736_5597# a_26036_4988.t49 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1188 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1189 a_24410_25128.t1 a_23436_16644.t46 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X1190 Vdd a_4288_11726# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1191 a_14832_12082.t0 a_14188_14050.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1192 a_22629_17217# Fvco.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1193 a_28478_5597# a_26036_4988.t50 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1194 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1195 a_50128_8156# a_54410_8156# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1196 a_28994_5597# a_26036_4988.t51 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1197 a_23160_10936.t1 a_14266_8900.t55 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1198 a_42574_15624# Fvco_By4_QPH_bar.t13 a_43010_16058# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1199 a_17685_3840.t3 vinit.t44 Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=1e+06u
X1200 a_27962_17218# a_26368_16652.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1201 a_25778_4988.t2 a_23414_5032.t46 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1202 a_54966_2992# a_49874_4150.t11 a_53308_2992# gnd sky130_fd_pr__nfet_01v8 ad=1.9575e+11p pd=1.64e+06u as=1.9575e+11p ps=1.64e+06u w=1.35e+06u l=8e+06u
X1203 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1204 a_25099_11445.t1 a_27762_11446.t47 a_17685_3840.t10 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1205 a_23160_10936.t0 a_14266_8900.t56 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1206 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1207 gnd gnd vinit.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1208 a_22972_23306.t3 vctrl a_17685_3840.t13 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1209 a_23156_5032.t1 a_14188_14050.t54 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1210 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1211 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1212 a_17685_3840.t12 vctrl a_22972_23306.t2 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1213 a_26589_17217# a_23436_16644.t47 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1214 a_8740_12844# Vso3b a_4226_11996# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1215 a_4314_11468# a_4226_11420# vout gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=1.0044e+12p ps=7.1e+06u w=3.24e+06u l=150000u
X1216 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1217 a_66154_26414# a_65077_26048# a_65992_26048# Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=5.88e+10p ps=700000u w=420000u l=150000u
X1218 a_27762_11446.t0 a_26368_16652.t52 a_17685_3840.t7 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1219 a_26589_17217# a_23436_16644.t48 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1220 a_38070_8852.t1 a_25099_11445.t53 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X1221 a_23178_16644# Fvco.t46 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1222 a_27962_17218# a_26368_16652.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1223 a_28478_5597# a_26036_4988.t52 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1224 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1225 gnd gnd vinit.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1226 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1227 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1228 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1229 a_22972_23306.t1 Vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X1230 a_51041_13108# Fvco_By4_QPH_bar.t14 a_50262_14152# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1231 a_25778_4988.t1 a_23414_5032.t47 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1232 a_26847_5596# a_23414_5032.t48 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1233 a_32948_24994.t0 a_27762_11446.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1234 a_28578_5014.t1 a_26036_4988.t53 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1235 a_63419_26414# RESET Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1236 a_28220_5597# a_26036_4988.t54 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1237 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1238 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1239 a_22629_5596# a_14188_14050.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1240 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1241 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1242 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1243 a_55602_11692# vbiasob.t4 a_51138_21494.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=2e+06u
X1244 a_23403_5596# a_14188_14050.t56 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1245 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1246 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1247 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1248 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1249 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1250 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1251 Vdd a_4226_11612# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1252 vbiasr.t1 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1253 Vdd Vdd vinit.t23 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1254 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1255 a_23661_17217# Fvco.t47 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1256 a_51041_13108# Fvco_By4_QPH_bar.t15 a_51276_14152# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.07143e+11p ps=1.67714e+06u w=1e+06u l=150000u
X1257 a_26847_5596# a_23414_5032.t49 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1258 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1259 a_26589_5596# a_23414_5032.t50 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1260 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1261 a_28220_5597# a_26036_4988.t55 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1262 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1263 Vdd a_64051_26022# a_64038_26414# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X1264 a_4314_11852# a_4226_11804# a_4314_11756# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X1265 a_26016_10878.t2 a_25099_11445.t54 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1266 gnd a_66178_25254# a_66742_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1267 a_26016_10878.t1 a_25099_11445.t55 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1268 a_28736_5597# a_26036_4988.t56 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1269 a_29510_5597# a_26036_4988.t57 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1270 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1271 aa vbiasbuffer.t4 a_50032_16080.t0 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=1e+06u
X1272 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1273 a_26847_11500# a_25099_11445.t56 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1274 a_51636_13108# Fvco_By4_QPH_bar.t16 a_50262_14152# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.07143e+11p ps=1.67714e+06u w=1e+06u l=150000u
X1275 vinit.t5 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1276 Vdd a_66003_25280# a_66178_25254# Vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X1277 a_8748_11692# Vso5b a_4226_11804# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1278 a_26073_11500# a_25099_11445.t57 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1279 gnd gnd vbiasr.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1280 Vdd Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1281 a_50262_14152# Fvco_By4_QPH.t16 a_51636_13108# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1282 a_23156_5032.t0 a_14188_14050.t57 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1283 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1284 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1285 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1286 CLK_BY_2_BAR.t1 a_64615_26048# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X1287 a_8744_9386# CLK_IN a_4226_11420# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1288 gnd a_17685_3840.t59 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1289 a_26589_5596# a_23414_5032.t51 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1290 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1291 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1292 a_26110_16652# a_23436_16644.t49 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1293 a_25299_17217# a_23436_16644.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1294 a_26073_11500# a_25099_11445.t58 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1295 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1296 a_65427_26048# a_64911_26048# a_65332_26048# gnd sky130_fd_pr__nfet_01v8 ad=5.94e+10p pd=690000u as=6.09231e+10p ps=687692u w=360000u l=150000u
X1297 Vdd a_64725_25280# a_64922_25280# Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1298 a_25299_17217# a_23436_16644.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1299 gnd a_17685_3840.t60 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1300 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1301 a_44752_16348.t2 bb a_42782_16060# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1302 a_25815_5596# a_23414_5032.t52 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1303 vinit.t4 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1304 a_27962_17218# a_26368_16652.t54 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1305 a_26331_5596# a_23414_5032.t53 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1306 gnd a_17685_3840.t61 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1307 a_28478_5597# a_26036_4988.t58 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1308 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1309 a_66178_25254# a_66003_25280# a_66357_25280# gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=6.405e+10p ps=725000u w=420000u l=150000u
X1310 gnd Vso8b a_8752_10532# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1311 a_29252_5597# a_26036_4988.t59 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1312 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1313 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1314 a_26073_17217# a_23436_16644.t52 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1315 a_27962_17218# a_26368_16652.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1316 a_25778_4988.t0 a_23414_5032.t54 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1317 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1318 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1319 a_47760_15642# a_43010_16058# a_33808_31746# Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.08286e+07u as=9.47286e+11p ps=7.07857e+06u w=5e+06u l=1e+06u
X1320 a_63529_26290# a_63311_26048# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.722e+11p pd=1.58e+06u as=1.81761e+11p ps=1.31123e+06u w=840000u l=150000u
X1321 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1322 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1323 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1324 a_23403_17217# Fvco.t48 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1325 a_4314_11948# a_4288_11918# a_4314_11852# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X1326 gnd a_17685_3840.t62 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1327 a_23178_16644# Fvco.t49 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1328 a_51532_4150.t2 a_49874_4150.t12 a_54966_3580# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.0035e+11p ps=5.12e+06u w=4.83e+06u l=8e+06u
X1329 a_77598_24640.t4 a_77572_23336.t0 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1330 gnd CLK_BY_2_BAR.t8 a_64725_25280# gnd sky130_fd_pr__nfet_01v8 ad=1.42392e+11p pd=1.0559e+06u as=8.775e+10p ps=920000u w=650000u l=150000u
X1331 a_23178_16644# Fvco.t50 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1332 a_25557_5596# a_23414_5032.t55 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1333 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1334 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1335 a_44752_16348.t0 aa a_42574_15624# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1336 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1337 a_26331_5596# a_23414_5032.t56 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1338 vinit.t22 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1339 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.416e+07u w=2.4e+07u
X1340 gnd Vso6b a_8748_11692# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1341 a_28994_11501# a_27762_11446.t49 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1342 a_26847_5596# a_23414_5032.t57 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1343 a_65332_26048# Fvco_By4_QPH.t17 Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=6.51e+10p pd=730000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1344 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1345 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1346 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1347 a_25815_11500# a_25099_11445.t59 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1348 a_28220_5597# a_26036_4988.t60 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1349 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1350 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1351 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1352 a_25815_11500# a_25099_11445.t60 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1353 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1354 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1355 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1356 a_8748_9956# Vso8b a_4288_11534# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1357 gnd a_17685_3840.t63 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1358 vinit.t3 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1359 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1360 a_25557_11500# a_25099_11445.t61 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1361 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1362 a_28994_11501# a_27762_11446.t50 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1363 a_25299_5596# a_23414_5032.t58 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1364 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1365 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1366 gnd gnd vinit.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1367 a_66178_25254# RESET Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1368 a_28994_11501# a_27762_11446.t51 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1369 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1370 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1371 Vdd a_4288_12110# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1372 a_25815_17217# a_23436_16644.t53 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1373 a_26589_5596# a_23414_5032.t59 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1374 a_28994_11501# a_27762_11446.t52 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1375 Vso8b a_30384_802.t3 Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1376 gnd a_66167_26022# a_66731_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1377 a_29510_11501# a_27762_11446.t53 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1378 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1379 a_24177_11500# a_14266_8900.t57 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1380 a_33808_31746# a_43010_16058# a_47760_15642# Vdd sky130_fd_pr__pfet_01v8_lvt ad=9.47286e+11p pd=7.07857e+06u as=1.45e+12p ps=1.08286e+07u w=5e+06u l=1e+06u
X1381 a.t0 a_77254_23336.t6 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1382 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1383 a_29510_11501# a_27762_11446.t54 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1384 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1385 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1386 a_28994_17218# a_26368_16652.t56 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1387 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1388 gnd a_17685_3840.t64 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1389 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1390 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1391 a_29252_11501# a_27762_11446.t55 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1392 a_42782_16060# Fvco_By4_QPH_bar.t17 a_42550_16062# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1393 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1394 gnd a_64051_26022# a_63985_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=7.20462e+10p ps=807692u w=420000u l=150000u
X1395 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1396 a_26110_16652# a_23436_16644.t54 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1397 a_50320_14126# Fvco_By4_QPH.t18 a_56602_11692# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X1398 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1399 a_29510_17218# a_26368_16652.t57 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1400 a_63985_26048# a_62795_26048# a_63876_26048# gnd sky130_fd_pr__nfet_01v8 ad=6.17538e+10p pd=692308u as=7.11e+10p ps=755000u w=360000u l=150000u
X1401 a_26110_16652# a_23436_16644.t55 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1402 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1403 vinit.t21 Vdd Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1404 a_28736_11501# a_27762_11446.t56 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1405 a_50262_14152# a_50320_14126# a_50511_16072.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X1406 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1407 a_66167_26022# a_65992_26048# a_66346_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=6.405e+10p ps=725000u w=420000u l=150000u
X1408 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1409 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1410 a_26073_17217# a_23436_16644.t56 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1411 a_51276_14152# a_51334_14126# a_33808_31746# gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=3.78571e+11p ps=2.99714e+06u w=2e+06u l=1e+06u
X1412 Vdd Vdd vinit.t20 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1413 a_26331_5596# a_23414_5032.t60 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1414 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1415 a_26073_17217# a_23436_16644.t57 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1416 Vdd a_4226_11804# vout Vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1417 a_29510_17218# a_26368_16652.t58 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1418 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1419 gnd gnd vinit.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1420 a_28736_11501# a_27762_11446.t57 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1421 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1422 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1423 a_65088_25280# a_64922_25280# Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.38484e+11p ps=999033u w=640000u l=150000u
X1424 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1425 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1426 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1427 a_28736_11501# a_27762_11446.t58 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1428 a_23919_5596# a_14188_14050.t58 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1429 a_50511_16072.t2 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1430 a_28736_11501# a_27762_11446.t59 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1431 gnd gnd vinit.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1432 a_23919_11500# a_14266_8900.t58 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1433 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1434 a_8736_14034# Vso1b a_4226_12188# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1435 a_65689_26048# a_65645_26290# a_65523_26048# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.50877e+11p ps=1.18462e+06u w=420000u l=150000u
X1436 a_28736_17218# a_26368_16652.t59 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1437 a_23145_11500# a_14266_8900.t59 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1438 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1439 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1440 a_23145_5596# a_14188_14050.t59 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1441 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1442 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1443 a_63876_26048# a_62961_26048# a_63529_26290# gnd sky130_fd_pr__nfet_01v8 ad=7.11e+10p pd=755000u as=7.1928e+10p ps=709200u w=360000u l=150000u
X1444 a_23145_11500# a_14266_8900.t60 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1445 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1446 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1447 a_65523_26048# a_65077_26048# a_65427_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.29323e+11p pd=1.01538e+06u as=5.94e+10p ps=690000u w=360000u l=150000u
X1448 gnd CLK_IN a_8748_9956# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1449 a_28220_11501# a_27762_11446.t60 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1450 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1451 a_22887_11500# a_14266_8900.t61 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1452 a_28220_11501# a_27762_11446.t61 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1453 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1454 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1455 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1456 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1457 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1458 a_23145_17217# Fvco.t4 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1459 a_77280_24640.t4 a_77254_23336.t2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1460 a_63216_26048# CLK_BY_2_BAR.t9 Vdd Vdd sky130_fd_pr__pfet_01v8_hvt ad=6.51e+10p pd=730000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1461 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1462 a_25815_17217# a_23436_16644.t58 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1463 Vdd Vdd vbiasr.t21 Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1464 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1465 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1466 a_28220_17218# a_26368_16652.t60 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1467 a_26589_17217# a_23436_16644.t59 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1468 a_26368_16652.t1 a_23436_16644.t60 a_17685_3840.t16 Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1469 a_25815_17217# a_23436_16644.t61 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1470 a_23145_5596# a_14188_14050.t60 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1471 a_8744_13422# Vso2b a_4288_12110# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1472 a_22887_5596# a_14188_14050.t61 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1473 aa Fvco_By4_QPH.t19 a_47760_15642# Vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.33143e+06u w=2e+06u l=150000u
X1474 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1475 a_8748_12270# Vso4b a_4288_11918# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1476 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1477 a_28994_17218# a_26368_16652.t61 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1478 a_28578_5014.t0 a_26036_4988.t61 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1479 Vdd a_34044_31208# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1480 Vdd a_9354_33563# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
C0 a_50262_14152# a_51636_13108# 2.25fF
C1 a_4226_12188# vout 2.67fF
C2 Vso3b Vdd 3.96fF
C3 a_55602_11692# a_56602_11692# 2.04fF
C4 a_9354_33563# a_33808_31746# 2.54fF
C5 Vdd a_9354_33563# 505.47fF
C6 a_51041_13108# a_51276_14152# 2.50fF
C7 a_47760_15642# a_47968_16078# 3.20fF
C8 Vdd CLK_BY_4_IPH 2.94fF
C9 a_55602_11692# a_51334_14126# 2.35fF
C10 CLK_IN vbiasr 2.24fF
C11 Vdd vinit 58.90fF
C12 Vso4b Vdd 3.85fF
C13 Fvco_By4_QPH Fvco_By4_QPH_bar 16.00fF
C14 Vso2b Vdd 3.24fF
C15 Vso6b Vdd 3.09fF
C16 a_47968_16078# aa 3.02fF
C17 a_42550_16062# a_42782_16060# 2.13fF
C18 Vdd CLK_BY_4_IPH_BAR 3.04fF
C19 vout Vdd 7.94fF
C20 a_47968_16078# bb 2.43fF
C21 a_42574_15624# a_43010_16058# 2.25fF
C22 vbiasr Vdd 50.30fF
C23 Fvco_By4_QPH RESET 2.21fF
C24 Vdd a_4226_11420# 2.26fF
C25 CLK_BY_4_IPH_BAR CLK_BY_4_IPH 2.04fF
C26 a_4288_12110# Vdd 2.60fF
C27 Vdd Fvco_By4_QPH_bar 2.21fF
C28 a_56602_11692# a_50320_14126# 2.53fF
C29 a_4226_11804# Vdd 2.43fF
C30 Vdd Vso7b 2.92fF
C31 a_4288_11918# Vdd 2.56fF
C32 a_50320_14126# a_51334_14126# 2.95fF
C33 a_50262_14152# a_51041_13108# 4.39fF
C34 Vso7b Vso8b 12.19fF
C35 a_4288_11726# Vdd 2.30fF
C36 Vso5b Vdd 5.20fF
C37 Vdd vbiasot 2.09fF
C38 Vso1b Vdd 3.70fF
C39 a_51041_13108# a_51636_13108# 4.40fF
C40 a_4226_11612# Vdd 2.37fF
C41 a_55602_11692# a_50320_14126# 2.15fF
C42 a_42550_16062# Vdd 5.00fF
C43 Vdd a_34044_31208# 504.99fF
C44 a_51636_13108# a_51276_14152# 2.56fF
C45 a_4288_11534# Vdd 2.42fF
C46 vctrl Vso1b 3.89fF
C47 a_47760_15642# aa 2.29fF
C48 a_42550_16062# a_42574_15624# 2.35fF
C49 a_4226_12188# Vdd 2.55fF
C50 Vso1b Vso2b 3.79fF
C51 a_47760_15642# bb 4.36fF
C52 a_42550_16062# a_43010_16058# 4.58fF
C53 a_42574_15624# a_42782_16060# 2.88fF
C54 CLK_IN Vdd 2.08fF
C55 a_42782_16060# a_43010_16058# 2.44fF
C56 vbiasob Vdd 3.11fF
C57 bb Fvco_By4_QPH_bar 2.30fF
C58 aa bb 2.62fF
C59 a_4226_11996# Vdd 2.88fF
C60 a_56602_11692# a_51334_14126# 2.10fF
C61 Vso4b CLK_IN 26.23fF
C62 a_51636_13108# a_56602_11692# 2.40fF
C63 a_33808_31746# a_51334_14126# 3.18fF
R0 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.n2 1158.04
R1 Fvco_By4_QPH_bar.t8 Fvco_By4_QPH_bar.t7 731.89
R2 Fvco_By4_QPH_bar.t3 Fvco_By4_QPH_bar.t12 719.978
R3 Fvco_By4_QPH_bar.t6 Fvco_By4_QPH_bar.t16 710.965
R4 Fvco_By4_QPH_bar.t5 Fvco_By4_QPH_bar.t17 710.965
R5 Fvco_By4_QPH_bar.t4 Fvco_By4_QPH_bar.t11 710.965
R6 Fvco_By4_QPH_bar.t16 Fvco_By4_QPH_bar.t15 579.889
R7 Fvco_By4_QPH_bar.t17 Fvco_By4_QPH_bar.t13 579.889
R8 Fvco_By4_QPH_bar.t11 Fvco_By4_QPH_bar.t10 579.889
R9 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.t5 570.03
R10 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.t4 563.963
R11 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t6 557.83
R12 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n0 458.189
R13 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.n5 435.858
R14 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t14 417.917
R15 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.t9 414.213
R16 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.t2 414.167
R17 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.t3 245.573
R18 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.t8 244.389
R19 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n7 188.615
R20 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n4 149.023
R21 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.n6 130.017
R22 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t0 69.215
R23 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n1 50.411
R24 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t1 39.949
R25 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.n3 1.452
R26 a_26368_16652.t24 a_26368_16652.t50 1273.78
R27 a_26368_16652.n3 a_26368_16652.t52 182.777
R28 a_26368_16652.n3 a_26368_16652.t1 127.728
R29 a_26368_16652.t52 a_26368_16652.t21 113.753
R30 a_26368_16652.t52 a_26368_16652.t27 113.753
R31 a_26368_16652.t52 a_26368_16652.t43 113.753
R32 a_26368_16652.t52 a_26368_16652.t59 113.753
R33 a_26368_16652.t52 a_26368_16652.t53 113.753
R34 a_26368_16652.t52 a_26368_16652.t3 113.753
R35 a_26368_16652.t52 a_26368_16652.t16 113.753
R36 a_26368_16652.t52 a_26368_16652.t32 113.753
R37 a_26368_16652.t39 a_26368_16652.t28 113.753
R38 a_26368_16652.t39 a_26368_16652.t42 113.753
R39 a_26368_16652.t39 a_26368_16652.t58 113.753
R40 a_26368_16652.t39 a_26368_16652.t12 113.753
R41 a_26368_16652.n0 a_26368_16652.t35 113.753
R42 a_26368_16652.n0 a_26368_16652.t48 113.753
R43 a_26368_16652.t39 a_26368_16652.t6 113.753
R44 a_26368_16652.t39 a_26368_16652.t61 113.753
R45 a_26368_16652.t39 a_26368_16652.t13 113.753
R46 a_26368_16652.t39 a_26368_16652.t29 113.753
R47 a_26368_16652.t39 a_26368_16652.t44 113.753
R48 a_26368_16652.n0 a_26368_16652.t22 113.753
R49 a_26368_16652.n0 a_26368_16652.t54 113.753
R50 a_26368_16652.n0 a_26368_16652.t8 113.753
R51 a_26368_16652.n0 a_26368_16652.t19 113.753
R52 a_26368_16652.t39 a_26368_16652.t37 113.753
R53 a_26368_16652.t39 a_26368_16652.t33 113.753
R54 a_26368_16652.t39 a_26368_16652.t46 113.753
R55 a_26368_16652.t39 a_26368_16652.t4 113.753
R56 a_26368_16652.t39 a_26368_16652.t17 113.753
R57 a_26368_16652.n0 a_26368_16652.t36 113.753
R58 a_26368_16652.n1 a_26368_16652.t49 113.753
R59 a_26368_16652.n1 a_26368_16652.t7 113.753
R60 a_26368_16652.t39 a_26368_16652.t2 113.753
R61 a_26368_16652.t39 a_26368_16652.t14 113.753
R62 a_26368_16652.t39 a_26368_16652.t30 113.753
R63 a_26368_16652.t39 a_26368_16652.t45 113.753
R64 a_26368_16652.n0 a_26368_16652.t23 113.753
R65 a_26368_16652.n0 a_26368_16652.t55 113.753
R66 a_26368_16652.n0 a_26368_16652.t9 113.753
R67 a_26368_16652.n2 a_26368_16652.t20 113.753
R68 a_26368_16652.n2 a_26368_16652.t38 113.753
R69 a_26368_16652.n2 a_26368_16652.t34 113.753
R70 a_26368_16652.n2 a_26368_16652.t47 113.753
R71 a_26368_16652.n2 a_26368_16652.t5 113.753
R72 a_26368_16652.n2 a_26368_16652.t18 113.753
R73 a_26368_16652.t52 a_26368_16652.t51 113.753
R74 a_26368_16652.t52 a_26368_16652.t60 113.753
R75 a_26368_16652.t52 a_26368_16652.t15 113.753
R76 a_26368_16652.t52 a_26368_16652.t31 113.753
R77 a_26368_16652.t39 a_26368_16652.t26 113.753
R78 a_26368_16652.t39 a_26368_16652.t41 113.753
R79 a_26368_16652.t39 a_26368_16652.t57 113.753
R80 a_26368_16652.t39 a_26368_16652.t11 113.753
R81 a_26368_16652.t52 a_26368_16652.t56 113.753
R82 a_26368_16652.t52 a_26368_16652.t10 113.753
R83 a_26368_16652.t52 a_26368_16652.t25 113.753
R84 a_26368_16652.t52 a_26368_16652.t40 113.753
R85 a_26368_16652.t0 a_26368_16652.n3 57.482
R86 a_26368_16652.t52 a_26368_16652.n0 5.834
R87 a_26368_16652.t39 a_26368_16652.n1 3.384
R88 a_26368_16652.t52 a_26368_16652.t24 3.018
R89 a_26368_16652.t39 a_26368_16652.n2 2.785
R90 a_26368_16652.t52 a_26368_16652.t39 2.574
R91 a_23414_5032.t2 a_23414_5032.t41 1273.78
R92 a_23414_5032.n4 a_23414_5032.t14 345.988
R93 a_23414_5032.n3 a_23414_5032.t5 113.753
R94 a_23414_5032.n3 a_23414_5032.t3 113.753
R95 a_23414_5032.n3 a_23414_5032.t15 113.753
R96 a_23414_5032.n2 a_23414_5032.t36 113.753
R97 a_23414_5032.n2 a_23414_5032.t33 113.753
R98 a_23414_5032.n2 a_23414_5032.t31 113.753
R99 a_23414_5032.n2 a_23414_5032.t30 113.753
R100 a_23414_5032.n0 a_23414_5032.t7 113.753
R101 a_23414_5032.n0 a_23414_5032.t39 113.753
R102 a_23414_5032.n0 a_23414_5032.t37 113.753
R103 a_23414_5032.n0 a_23414_5032.t34 113.753
R104 a_23414_5032.n0 a_23414_5032.t45 113.753
R105 a_23414_5032.t14 a_23414_5032.t11 113.753
R106 a_23414_5032.t14 a_23414_5032.t8 113.753
R107 a_23414_5032.t14 a_23414_5032.t6 113.753
R108 a_23414_5032.t14 a_23414_5032.t4 113.753
R109 a_23414_5032.n0 a_23414_5032.t21 113.753
R110 a_23414_5032.n0 a_23414_5032.t17 113.753
R111 a_23414_5032.n1 a_23414_5032.t35 113.753
R112 a_23414_5032.n1 a_23414_5032.t56 113.753
R113 a_23414_5032.n1 a_23414_5032.t51 113.753
R114 a_23414_5032.n1 a_23414_5032.t49 113.753
R115 a_23414_5032.n1 a_23414_5032.t47 113.753
R116 a_23414_5032.n0 a_23414_5032.t24 113.753
R117 a_23414_5032.n0 a_23414_5032.t58 113.753
R118 a_23414_5032.n0 a_23414_5032.t55 113.753
R119 a_23414_5032.n0 a_23414_5032.t52 113.753
R120 a_23414_5032.t14 a_23414_5032.t9 113.753
R121 a_23414_5032.t14 a_23414_5032.t28 113.753
R122 a_23414_5032.t14 a_23414_5032.t25 113.753
R123 a_23414_5032.t14 a_23414_5032.t23 113.753
R124 a_23414_5032.t14 a_23414_5032.t20 113.753
R125 a_23414_5032.n0 a_23414_5032.t27 113.753
R126 a_23414_5032.t14 a_23414_5032.t26 113.753
R127 a_23414_5032.t14 a_23414_5032.t42 113.753
R128 a_23414_5032.t14 a_23414_5032.t60 113.753
R129 a_23414_5032.t14 a_23414_5032.t59 113.753
R130 a_23414_5032.t14 a_23414_5032.t57 113.753
R131 a_23414_5032.t14 a_23414_5032.t54 113.753
R132 a_23414_5032.n0 a_23414_5032.t29 113.753
R133 a_23414_5032.n0 a_23414_5032.t13 113.753
R134 a_23414_5032.n0 a_23414_5032.t12 113.753
R135 a_23414_5032.t14 a_23414_5032.t10 113.753
R136 a_23414_5032.t14 a_23414_5032.t19 113.753
R137 a_23414_5032.t14 a_23414_5032.t44 113.753
R138 a_23414_5032.t14 a_23414_5032.t43 113.753
R139 a_23414_5032.t14 a_23414_5032.t40 113.753
R140 a_23414_5032.t14 a_23414_5032.t38 113.753
R141 a_23414_5032.n0 a_23414_5032.t22 113.753
R142 a_23414_5032.n0 a_23414_5032.t18 113.753
R143 a_23414_5032.n0 a_23414_5032.t16 113.753
R144 a_23414_5032.t14 a_23414_5032.t32 113.753
R145 a_23414_5032.t14 a_23414_5032.t53 113.753
R146 a_23414_5032.t14 a_23414_5032.t50 113.753
R147 a_23414_5032.t14 a_23414_5032.t48 113.753
R148 a_23414_5032.t14 a_23414_5032.t46 113.753
R149 a_23414_5032.t0 a_23414_5032.n5 82.513
R150 a_23414_5032.n4 a_23414_5032.t1 28.697
R151 a_23414_5032.t14 a_23414_5032.n0 4.31
R152 a_23414_5032.n5 a_23414_5032.n4 3.507
R153 a_23414_5032.n0 a_23414_5032.n3 3.224
R154 a_23414_5032.t14 a_23414_5032.n1 2.869
R155 a_23414_5032.t14 a_23414_5032.n2 2.708
R156 a_23414_5032.n5 a_23414_5032.t2 2.634
R157 a_26690_784.n1 a_26690_784.t2 434.481
R158 a_26690_784.n0 a_26690_784.t3 217.163
R159 a_26690_784.t1 a_26690_784.n1 52.152
R160 a_26690_784.n0 a_26690_784.t0 3.106
R161 a_26690_784.n1 a_26690_784.n0 0.879
R162 a_14188_14050.t12 a_14188_14050.t53 1273.78
R163 a_14188_14050.n3 a_14188_14050.t31 161.992
R164 a_14188_14050.t39 a_14188_14050.t40 113.753
R165 a_14188_14050.t39 a_14188_14050.t50 113.753
R166 a_14188_14050.t39 a_14188_14050.t47 113.753
R167 a_14188_14050.t39 a_14188_14050.t11 113.753
R168 a_14188_14050.n0 a_14188_14050.t23 113.753
R169 a_14188_14050.n0 a_14188_14050.t6 113.753
R170 a_14188_14050.n0 a_14188_14050.t19 113.753
R171 a_14188_14050.n0 a_14188_14050.t41 113.753
R172 a_14188_14050.t39 a_14188_14050.t55 113.753
R173 a_14188_14050.t39 a_14188_14050.t9 113.753
R174 a_14188_14050.t39 a_14188_14050.t8 113.753
R175 a_14188_14050.t39 a_14188_14050.t26 113.753
R176 a_14188_14050.n0 a_14188_14050.t42 113.753
R177 a_14188_14050.n0 a_14188_14050.t24 113.753
R178 a_14188_14050.n0 a_14188_14050.t38 113.753
R179 a_14188_14050.n0 a_14188_14050.t57 113.753
R180 a_14188_14050.t31 a_14188_14050.t21 113.753
R181 a_14188_14050.t31 a_14188_14050.t36 113.753
R182 a_14188_14050.t31 a_14188_14050.t33 113.753
R183 a_14188_14050.t31 a_14188_14050.t56 113.753
R184 a_14188_14050.n0 a_14188_14050.t10 113.753
R185 a_14188_14050.n0 a_14188_14050.t51 113.753
R186 a_14188_14050.n0 a_14188_14050.t5 113.753
R187 a_14188_14050.n0 a_14188_14050.t25 113.753
R188 a_14188_14050.t31 a_14188_14050.t49 113.753
R189 a_14188_14050.t31 a_14188_14050.t4 113.753
R190 a_14188_14050.t31 a_14188_14050.t60 113.753
R191 a_14188_14050.t31 a_14188_14050.t22 113.753
R192 a_14188_14050.n1 a_14188_14050.t37 113.753
R193 a_14188_14050.n1 a_14188_14050.t18 113.753
R194 a_14188_14050.n1 a_14188_14050.t30 113.753
R195 a_14188_14050.n1 a_14188_14050.t54 113.753
R196 a_14188_14050.n2 a_14188_14050.t3 113.753
R197 a_14188_14050.n2 a_14188_14050.t16 113.753
R198 a_14188_14050.n2 a_14188_14050.t14 113.753
R199 a_14188_14050.n2 a_14188_14050.t35 113.753
R200 a_14188_14050.n0 a_14188_14050.t48 113.753
R201 a_14188_14050.n0 a_14188_14050.t29 113.753
R202 a_14188_14050.n0 a_14188_14050.t45 113.753
R203 a_14188_14050.n0 a_14188_14050.t7 113.753
R204 a_14188_14050.t31 a_14188_14050.t46 113.753
R205 a_14188_14050.t31 a_14188_14050.t61 113.753
R206 a_14188_14050.t31 a_14188_14050.t59 113.753
R207 a_14188_14050.t31 a_14188_14050.t20 113.753
R208 a_14188_14050.t31 a_14188_14050.t28 113.753
R209 a_14188_14050.t31 a_14188_14050.t44 113.753
R210 a_14188_14050.t31 a_14188_14050.t43 113.753
R211 a_14188_14050.t31 a_14188_14050.t2 113.753
R212 a_14188_14050.n0 a_14188_14050.t15 113.753
R213 a_14188_14050.n0 a_14188_14050.t58 113.753
R214 a_14188_14050.n0 a_14188_14050.t13 113.753
R215 a_14188_14050.n0 a_14188_14050.t32 113.753
R216 a_14188_14050.t31 a_14188_14050.t34 113.753
R217 a_14188_14050.t31 a_14188_14050.t17 113.753
R218 a_14188_14050.t31 a_14188_14050.t27 113.753
R219 a_14188_14050.n0 a_14188_14050.t52 113.753
R220 a_14188_14050.t1 a_14188_14050.n4 57.821
R221 a_14188_14050.n3 a_14188_14050.t0 47.07
R222 a_14188_14050.n4 a_14188_14050.t12 6.878
R223 a_14188_14050.n4 a_14188_14050.n3 3.96
R224 a_14188_14050.t31 a_14188_14050.t39 3.88
R225 a_14188_14050.t31 a_14188_14050.n0 3.25
R226 a_14188_14050.n0 a_14188_14050.n1 2.856
R227 a_14188_14050.t31 a_14188_14050.n2 2.454
R228 a_49874_4150.n0 a_49874_4150.t12 19.742
R229 a_49874_4150.n0 a_49874_4150.t6 18.733
R230 a_49874_4150.t0 a_49874_4150.n1 18.498
R231 a_49874_4150.n3 a_49874_4150.t3 17.928
R232 a_49874_4150.n0 a_49874_4150.t9 16.208
R233 a_49874_4150.n1 a_49874_4150.t2 15.946
R234 a_49874_4150.n2 a_49874_4150.t5 9.424
R235 a_49874_4150.n2 a_49874_4150.t8 8.34
R236 a_49874_4150.n2 a_49874_4150.t11 5.724
R237 a_49874_4150.n1 a_49874_4150.t1 5.514
R238 a_49874_4150.n0 a_49874_4150.t4 5.514
R239 a_49874_4150.n3 a_49874_4150.t7 5.512
R240 a_49874_4150.n1 a_49874_4150.n0 4.479
R241 a_49874_4150.n4 a_49874_4150.n3 4.094
R242 a_49874_4150.n4 a_49874_4150.t10 3.856
R243 a_49874_4150.n0 a_49874_4150.n4 3.301
R244 a_49874_4150.n0 a_49874_4150.n2 2.294
R245 Fvco_By4_QPH.t10 Fvco_By4_QPH.t19 731.89
R246 Fvco_By4_QPH.t14 Fvco_By4_QPH.t6 731.89
R247 Fvco_By4_QPH.t3 Fvco_By4_QPH.t13 731.89
R248 Fvco_By4_QPH.t5 Fvco_By4_QPH.t16 718.506
R249 Fvco_By4_QPH.t11 Fvco_By4_QPH.t15 710.965
R250 Fvco_By4_QPH.t7 Fvco_By4_QPH.t14 622.637
R251 Fvco_By4_QPH.n8 Fvco_By4_QPH.n7 617.524
R252 Fvco_By4_QPH.n4 Fvco_By4_QPH.n3 580.872
R253 Fvco_By4_QPH.t15 Fvco_By4_QPH.t2 579.889
R254 Fvco_By4_QPH.n3 Fvco_By4_QPH.t12 491.229
R255 Fvco_By4_QPH.n4 Fvco_By4_QPH.t4 489.182
R256 Fvco_By4_QPH.n9 Fvco_By4_QPH.t11 418.965
R257 Fvco_By4_QPH.n8 Fvco_By4_QPH.t18 414.13
R258 Fvco_By4_QPH.n5 Fvco_By4_QPH.t9 349.273
R259 Fvco_By4_QPH.n2 Fvco_By4_QPH.t8 333.651
R260 Fvco_By4_QPH.n6 Fvco_By4_QPH.t3 317.894
R261 Fvco_By4_QPH.n2 Fvco_By4_QPH.t17 297.233
R262 Fvco_By4_QPH.n6 Fvco_By4_QPH.t5 291.323
R263 Fvco_By4_QPH.n5 Fvco_By4_QPH.t10 252.624
R264 Fvco_By4_QPH.n3 Fvco_By4_QPH.t7 227.612
R265 Fvco_By4_QPH.t9 Fvco_By4_QPH.n4 227.612
R266 Fvco_By4_QPH.n7 Fvco_By4_QPH.n5 198.896
R267 Fvco_By4_QPH.n9 Fvco_By4_QPH.n8 152.778
R268 Fvco_By4_QPH.n0 Fvco_By4_QPH.t1 92.046
R269 Fvco_By4_QPH.n1 Fvco_By4_QPH.n2 70.221
R270 Fvco_By4_QPH.n0 Fvco_By4_QPH.t0 61.427
R271 Fvco_By4_QPH Fvco_By4_QPH.n9 38.508
R272 Fvco_By4_QPH.n7 Fvco_By4_QPH.n6 31.687
R273 Fvco_By4_QPH Fvco_By4_QPH.n1 10.972
R274 Fvco_By4_QPH.n1 Fvco_By4_QPH.n0 0.154
R275 vbiasr.n16 vbiasr.t20 11.76
R276 vbiasr.n27 vbiasr.t29 7.425
R277 vbiasr.n16 vbiasr.t35 7.425
R278 vbiasr.n25 vbiasr.t28 5.713
R279 vbiasr.n25 vbiasr.t36 5.713
R280 vbiasr.n8 vbiasr.t21 5.713
R281 vbiasr.n8 vbiasr.t40 5.713
R282 vbiasr.n9 vbiasr.t26 5.713
R283 vbiasr.n9 vbiasr.t24 5.713
R284 vbiasr.n10 vbiasr.t23 5.713
R285 vbiasr.n10 vbiasr.t30 5.713
R286 vbiasr.n12 vbiasr.t34 5.713
R287 vbiasr.n12 vbiasr.t33 5.713
R288 vbiasr.n13 vbiasr.t27 5.713
R289 vbiasr.n13 vbiasr.t25 5.713
R290 vbiasr.n14 vbiasr.t31 5.713
R291 vbiasr.n14 vbiasr.t22 5.713
R292 vbiasr.n15 vbiasr.t32 5.713
R293 vbiasr.n15 vbiasr.t37 5.713
R294 vbiasr.n11 vbiasr.t39 5.713
R295 vbiasr.n11 vbiasr.t38 5.713
R296 vbiasr.n39 vbiasr.t1 5.244
R297 vbiasr.n28 vbiasr.t7 5.244
R298 vbiasr.n0 vbiasr.t13 3.48
R299 vbiasr.n0 vbiasr.t8 3.48
R300 vbiasr.n1 vbiasr.t5 3.48
R301 vbiasr.n1 vbiasr.t11 3.48
R302 vbiasr.n2 vbiasr.t10 3.48
R303 vbiasr.n2 vbiasr.t12 3.48
R304 vbiasr.n3 vbiasr.t17 3.48
R305 vbiasr.n3 vbiasr.t16 3.48
R306 vbiasr.n4 vbiasr.t0 3.48
R307 vbiasr.n4 vbiasr.t9 3.48
R308 vbiasr.n5 vbiasr.t6 3.48
R309 vbiasr.n5 vbiasr.t4 3.48
R310 vbiasr.n6 vbiasr.t3 3.48
R311 vbiasr.n6 vbiasr.t19 3.48
R312 vbiasr.n7 vbiasr.t18 3.48
R313 vbiasr.n7 vbiasr.t15 3.48
R314 vbiasr.n29 vbiasr.t14 3.48
R315 vbiasr.n29 vbiasr.t2 3.48
R316 vbiasr.n35 vbiasr.n3 1.766
R317 vbiasr.n38 vbiasr.n0 1.766
R318 vbiasr.n32 vbiasr.n6 1.766
R319 vbiasr.n31 vbiasr.n7 1.764
R320 vbiasr.n34 vbiasr.n4 1.762
R321 vbiasr.n36 vbiasr.n2 1.761
R322 vbiasr.n33 vbiasr.n5 1.758
R323 vbiasr.n37 vbiasr.n1 1.758
R324 vbiasr.n30 vbiasr.n29 1.754
R325 vbiasr.n20 vbiasr.n12 1.714
R326 vbiasr.n17 vbiasr.n15 1.714
R327 vbiasr.n23 vbiasr.n9 1.714
R328 vbiasr.n24 vbiasr.n8 1.712
R329 vbiasr.n21 vbiasr.n11 1.71
R330 vbiasr.n19 vbiasr.n13 1.709
R331 vbiasr.n22 vbiasr.n10 1.706
R332 vbiasr.n18 vbiasr.n14 1.706
R333 vbiasr.n26 vbiasr.n25 1.702
R334 vbiasr.n28 vbiasr.n27 0.292
R335 vbiasr vbiasr.n39 0.152
R336 vbiasr.n22 vbiasr.n21 0.031
R337 vbiasr.n34 vbiasr.n33 0.031
R338 vbiasr.n19 vbiasr.n18 0.031
R339 vbiasr.n37 vbiasr.n36 0.031
R340 vbiasr.n31 vbiasr.n30 0.031
R341 vbiasr.n26 vbiasr.n24 0.031
R342 vbiasr.n30 vbiasr.n28 0.031
R343 vbiasr.n27 vbiasr.n26 0.031
R344 vbiasr.n38 vbiasr.n37 0.03
R345 vbiasr.n18 vbiasr.n17 0.03
R346 vbiasr.n39 vbiasr.n38 0.03
R347 vbiasr.n17 vbiasr.n16 0.03
R348 vbiasr.n24 vbiasr.n23 0.03
R349 vbiasr.n32 vbiasr.n31 0.03
R350 vbiasr.n21 vbiasr.n20 0.03
R351 vbiasr.n35 vbiasr.n34 0.03
R352 vbiasr.n20 vbiasr.n19 0.03
R353 vbiasr.n36 vbiasr.n35 0.03
R354 vbiasr.n33 vbiasr.n32 0.03
R355 vbiasr.n23 vbiasr.n22 0.03
R356 a_26036_4988.t16 a_26036_4988.t22 1273.78
R357 a_26036_4988.n0 a_26036_4988.t44 415.476
R358 a_26036_4988.t44 a_26036_4988.t37 113.753
R359 a_26036_4988.t44 a_26036_4988.t34 113.753
R360 a_26036_4988.t44 a_26036_4988.t32 113.753
R361 a_26036_4988.t20 a_26036_4988.t46 113.753
R362 a_26036_4988.t20 a_26036_4988.t7 113.753
R363 a_26036_4988.t20 a_26036_4988.t4 113.753
R364 a_26036_4988.t20 a_26036_4988.t61 113.753
R365 a_26036_4988.t44 a_26036_4988.t14 113.753
R366 a_26036_4988.t44 a_26036_4988.t47 113.753
R367 a_26036_4988.t44 a_26036_4988.t10 113.753
R368 a_26036_4988.t44 a_26036_4988.t6 113.753
R369 a_26036_4988.t44 a_26036_4988.t3 113.753
R370 a_26036_4988.t20 a_26036_4988.t15 113.753
R371 a_26036_4988.t20 a_26036_4988.t41 113.753
R372 a_26036_4988.t20 a_26036_4988.t38 113.753
R373 a_26036_4988.t20 a_26036_4988.t35 113.753
R374 a_26036_4988.n1 a_26036_4988.t55 113.753
R375 a_26036_4988.n1 a_26036_4988.t52 113.753
R376 a_26036_4988.t20 a_26036_4988.t49 113.753
R377 a_26036_4988.t20 a_26036_4988.t5 113.753
R378 a_26036_4988.t20 a_26036_4988.t27 113.753
R379 a_26036_4988.t20 a_26036_4988.t25 113.753
R380 a_26036_4988.t20 a_26036_4988.t18 113.753
R381 a_26036_4988.n1 a_26036_4988.t36 113.753
R382 a_26036_4988.n1 a_26036_4988.t8 113.753
R383 a_26036_4988.n1 a_26036_4988.t29 113.753
R384 a_26036_4988.n1 a_26036_4988.t26 113.753
R385 a_26036_4988.t20 a_26036_4988.t23 113.753
R386 a_26036_4988.t20 a_26036_4988.t39 113.753
R387 a_26036_4988.t20 a_26036_4988.t59 113.753
R388 a_26036_4988.t20 a_26036_4988.t57 113.753
R389 a_26036_4988.t20 a_26036_4988.t53 113.753
R390 a_26036_4988.n1 a_26036_4988.t60 113.753
R391 a_26036_4988.t20 a_26036_4988.t58 113.753
R392 a_26036_4988.t20 a_26036_4988.t56 113.753
R393 a_26036_4988.t20 a_26036_4988.t11 113.753
R394 a_26036_4988.t20 a_26036_4988.t31 113.753
R395 a_26036_4988.t20 a_26036_4988.t30 113.753
R396 a_26036_4988.t20 a_26036_4988.t28 113.753
R397 a_26036_4988.n1 a_26036_4988.t42 113.753
R398 a_26036_4988.n1 a_26036_4988.t19 113.753
R399 a_26036_4988.n1 a_26036_4988.t45 113.753
R400 a_26036_4988.n2 a_26036_4988.t43 113.753
R401 a_26036_4988.n2 a_26036_4988.t40 113.753
R402 a_26036_4988.n2 a_26036_4988.t51 113.753
R403 a_26036_4988.n2 a_26036_4988.t13 113.753
R404 a_26036_4988.n2 a_26036_4988.t12 113.753
R405 a_26036_4988.n2 a_26036_4988.t9 113.753
R406 a_26036_4988.t44 a_26036_4988.t33 113.753
R407 a_26036_4988.t44 a_26036_4988.t54 113.753
R408 a_26036_4988.t44 a_26036_4988.t50 113.753
R409 a_26036_4988.t44 a_26036_4988.t48 113.753
R410 a_26036_4988.t44 a_26036_4988.t2 113.753
R411 a_26036_4988.t44 a_26036_4988.t24 113.753
R412 a_26036_4988.t44 a_26036_4988.t21 113.753
R413 a_26036_4988.t44 a_26036_4988.t17 113.753
R414 a_26036_4988.t1 a_26036_4988.n0 81.094
R415 a_26036_4988.n0 a_26036_4988.t0 28.577
R416 a_26036_4988.t44 a_26036_4988.n1 6.49
R417 a_26036_4988.n0 a_26036_4988.t16 5.37
R418 a_26036_4988.t20 a_26036_4988.n2 4.699
R419 a_26036_4988.t44 a_26036_4988.t20 2.967
R420 CLK_BY_4_IPH.n0 CLK_BY_4_IPH.t6 440.519
R421 CLK_BY_4_IPH.n0 CLK_BY_4_IPH.t5 402.739
R422 CLK_BY_4_IPH.n2 CLK_BY_4_IPH.t4 227.612
R423 CLK_BY_4_IPH.n1 CLK_BY_4_IPH.t3 227.612
R424 CLK_BY_4_IPH.n1 CLK_BY_4_IPH.n0 183.872
R425 CLK_BY_4_IPH.n3 CLK_BY_4_IPH.n2 179.1
R426 CLK_BY_4_IPH CLK_BY_4_IPH.t1 57.015
R427 CLK_BY_4_IPH.n2 CLK_BY_4_IPH.n1 45.046
R428 CLK_BY_4_IPH.n4 CLK_BY_4_IPH.t2 40.318
R429 CLK_BY_4_IPH.n3 CLK_BY_4_IPH.t0 15.901
R430 CLK_BY_4_IPH CLK_BY_4_IPH.n4 11.83
R431 CLK_BY_4_IPH.n4 CLK_BY_4_IPH.n3 0.329
R432 a_25099_11445.t53 a_25099_11445.t41 1273.78
R433 a_25099_11445.n3 a_25099_11445.t40 218.051
R434 a_25099_11445.t40 a_25099_11445.t49 113.753
R435 a_25099_11445.t40 a_25099_11445.t8 113.753
R436 a_25099_11445.t40 a_25099_11445.t29 113.753
R437 a_25099_11445.t40 a_25099_11445.t21 113.753
R438 a_25099_11445.t40 a_25099_11445.t42 113.753
R439 a_25099_11445.t40 a_25099_11445.t59 113.753
R440 a_25099_11445.t40 a_25099_11445.t57 113.753
R441 a_25099_11445.n2 a_25099_11445.t6 113.753
R442 a_25099_11445.n2 a_25099_11445.t16 113.753
R443 a_25099_11445.n2 a_25099_11445.t37 113.753
R444 a_25099_11445.n2 a_25099_11445.t54 113.753
R445 a_25099_11445.t40 a_25099_11445.t19 113.753
R446 a_25099_11445.n0 a_25099_11445.t51 113.753
R447 a_25099_11445.n0 a_25099_11445.t10 113.753
R448 a_25099_11445.n0 a_25099_11445.t31 113.753
R449 a_25099_11445.n1 a_25099_11445.t26 113.753
R450 a_25099_11445.n1 a_25099_11445.t35 113.753
R451 a_25099_11445.n1 a_25099_11445.t47 113.753
R452 a_25099_11445.n1 a_25099_11445.t4 113.753
R453 a_25099_11445.n1 a_25099_11445.t23 113.753
R454 a_25099_11445.n0 a_25099_11445.t43 113.753
R455 a_25099_11445.n0 a_25099_11445.t60 113.753
R456 a_25099_11445.t15 a_25099_11445.t58 113.753
R457 a_25099_11445.t15 a_25099_11445.t7 113.753
R458 a_25099_11445.t15 a_25099_11445.t17 113.753
R459 a_25099_11445.t15 a_25099_11445.t38 113.753
R460 a_25099_11445.t15 a_25099_11445.t55 113.753
R461 a_25099_11445.n0 a_25099_11445.t20 113.753
R462 a_25099_11445.n0 a_25099_11445.t52 113.753
R463 a_25099_11445.n0 a_25099_11445.t11 113.753
R464 a_25099_11445.t15 a_25099_11445.t32 113.753
R465 a_25099_11445.t15 a_25099_11445.t27 113.753
R466 a_25099_11445.t15 a_25099_11445.t36 113.753
R467 a_25099_11445.t15 a_25099_11445.t48 113.753
R468 a_25099_11445.t15 a_25099_11445.t5 113.753
R469 a_25099_11445.t15 a_25099_11445.t24 113.753
R470 a_25099_11445.t15 a_25099_11445.t39 113.753
R471 a_25099_11445.t15 a_25099_11445.t56 113.753
R472 a_25099_11445.t15 a_25099_11445.t12 113.753
R473 a_25099_11445.n0 a_25099_11445.t44 113.753
R474 a_25099_11445.n0 a_25099_11445.t61 113.753
R475 a_25099_11445.t15 a_25099_11445.t14 113.753
R476 a_25099_11445.t15 a_25099_11445.t13 113.753
R477 a_25099_11445.t15 a_25099_11445.t28 113.753
R478 a_25099_11445.t40 a_25099_11445.t50 113.753
R479 a_25099_11445.t40 a_25099_11445.t9 113.753
R480 a_25099_11445.t40 a_25099_11445.t30 113.753
R481 a_25099_11445.t40 a_25099_11445.t25 113.753
R482 a_25099_11445.t15 a_25099_11445.t34 113.753
R483 a_25099_11445.t15 a_25099_11445.t46 113.753
R484 a_25099_11445.t15 a_25099_11445.t3 113.753
R485 a_25099_11445.t15 a_25099_11445.t22 113.753
R486 a_25099_11445.t40 a_25099_11445.t33 113.753
R487 a_25099_11445.t40 a_25099_11445.t45 113.753
R488 a_25099_11445.t40 a_25099_11445.t2 113.753
R489 a_25099_11445.t40 a_25099_11445.t18 113.753
R490 a_25099_11445.t0 a_25099_11445.n4 56.779
R491 a_25099_11445.n3 a_25099_11445.t1 28.581
R492 a_25099_11445.t40 a_25099_11445.n0 5.834
R493 a_25099_11445.n4 a_25099_11445.t53 4.799
R494 a_25099_11445.n4 a_25099_11445.n3 3.709
R495 a_25099_11445.t15 a_25099_11445.n1 2.869
R496 a_25099_11445.t40 a_25099_11445.t15 2.816
R497 a_25099_11445.t15 a_25099_11445.n2 2.586
R498 a_17685_3840.n28 a_17685_3840.n27 660.793
R499 a_17685_3840.n56 a_17685_3840.n55 649.743
R500 a_17685_3840.n61 a_17685_3840.n60 574.593
R501 a_17685_3840.n29 a_17685_3840.n28 416.406
R502 a_17685_3840.n62 a_17685_3840.n61 415.789
R503 a_17685_3840.n58 a_17685_3840.n57 271.45
R504 a_17685_3840.n60 a_17685_3840.n59 262.496
R505 a_17685_3840.n28 a_17685_3840.n26 198.935
R506 a_17685_3840.n60 a_17685_3840.t11 197.212
R507 a_17685_3840.n59 a_17685_3840.t9 185.816
R508 a_17685_3840.n27 a_17685_3840.t15 176.327
R509 a_17685_3840.n58 a_17685_3840.t4 173.989
R510 a_17685_3840.n26 a_17685_3840.t10 154.605
R511 a_17685_3840.n57 a_17685_3840.t6 151.674
R512 a_17685_3840.n63 a_17685_3840.t5 118.032
R513 a_17685_3840.n61 a_17685_3840.n58 107.97
R514 a_17685_3840.n30 a_17685_3840.n29 104.297
R515 a_17685_3840.n64 a_17685_3840.n63 103.649
R516 a_17685_3840.n32 a_17685_3840.n1 100.878
R517 a_17685_3840.n65 a_17685_3840.n64 83.404
R518 a_17685_3840.n65 a_17685_3840.t16 81.437
R519 a_17685_3840.n30 a_17685_3840.t7 69.653
R520 a_17685_3840.n31 a_17685_3840.t1 68.683
R521 a_17685_3840.n64 a_17685_3840.n0 66.545
R522 a_17685_3840.n63 a_17685_3840.n62 47.861
R523 a_17685_3840.n25 a_17685_3840.n24 45.936
R524 a_17685_3840.n31 a_17685_3840.n30 45.7
R525 a_17685_3840.n29 a_17685_3840.n25 41.108
R526 a_17685_3840.n62 a_17685_3840.n56 41.07
R527 a_17685_3840.n67 a_17685_3840.n66 40.119
R528 a_17685_3840.n0 a_17685_3840.t13 29.277
R529 a_17685_3840.n0 a_17685_3840.t12 28.576
R530 a_17685_3840.n0 a_17685_3840.t14 28.565
R531 a_17685_3840.n1 a_17685_3840.t2 28.565
R532 a_17685_3840.n1 a_17685_3840.t8 28.565
R533 a_17685_3840.t0 a_17685_3840.n67 28.565
R534 a_17685_3840.n67 a_17685_3840.t3 28.565
R535 a_17685_3840.n55 a_17685_3840.n43 24.999
R536 a_17685_3840.n66 a_17685_3840.n65 24.605
R537 a_17685_3840.n24 a_17685_3840.n12 24.399
R538 a_17685_3840.n33 a_17685_3840.t50 23.529
R539 a_17685_3840.n2 a_17685_3840.t43 23.485
R540 a_17685_3840.n13 a_17685_3840.t35 23.474
R541 a_17685_3840.n44 a_17685_3840.t59 23.456
R542 a_17685_3840.n66 a_17685_3840.n32 20.217
R543 a_17685_3840.n32 a_17685_3840.n31 19.791
R544 a_17685_3840.n43 a_17685_3840.t39 15.401
R545 a_17685_3840.n12 a_17685_3840.t54 15.374
R546 a_17685_3840.n54 a_17685_3840.t26 15.341
R547 a_17685_3840.n23 a_17685_3840.t27 15.334
R548 a_17685_3840.n24 a_17685_3840.n23 12.228
R549 a_17685_3840.n55 a_17685_3840.n54 11.433
R550 a_17685_3840.n42 a_17685_3840.n41 10.674
R551 a_17685_3840.n41 a_17685_3840.n40 10.674
R552 a_17685_3840.n40 a_17685_3840.n39 10.674
R553 a_17685_3840.n39 a_17685_3840.n38 10.674
R554 a_17685_3840.n38 a_17685_3840.n37 10.674
R555 a_17685_3840.n37 a_17685_3840.n36 10.674
R556 a_17685_3840.n36 a_17685_3840.n35 10.674
R557 a_17685_3840.n35 a_17685_3840.n34 10.674
R558 a_17685_3840.n34 a_17685_3840.n33 10.674
R559 a_17685_3840.n22 a_17685_3840.n21 10.655
R560 a_17685_3840.n21 a_17685_3840.n20 10.655
R561 a_17685_3840.n20 a_17685_3840.n19 10.655
R562 a_17685_3840.n19 a_17685_3840.n18 10.655
R563 a_17685_3840.n18 a_17685_3840.n17 10.655
R564 a_17685_3840.n17 a_17685_3840.n16 10.655
R565 a_17685_3840.n16 a_17685_3840.n15 10.655
R566 a_17685_3840.n15 a_17685_3840.n14 10.655
R567 a_17685_3840.n14 a_17685_3840.n13 10.655
R568 a_17685_3840.n11 a_17685_3840.n10 10.637
R569 a_17685_3840.n10 a_17685_3840.n9 10.637
R570 a_17685_3840.n9 a_17685_3840.n8 10.637
R571 a_17685_3840.n8 a_17685_3840.n7 10.637
R572 a_17685_3840.n7 a_17685_3840.n6 10.637
R573 a_17685_3840.n6 a_17685_3840.n5 10.637
R574 a_17685_3840.n5 a_17685_3840.n4 10.637
R575 a_17685_3840.n4 a_17685_3840.n3 10.637
R576 a_17685_3840.n3 a_17685_3840.n2 10.637
R577 a_17685_3840.n53 a_17685_3840.n52 10.625
R578 a_17685_3840.n52 a_17685_3840.n51 10.625
R579 a_17685_3840.n51 a_17685_3840.n50 10.625
R580 a_17685_3840.n50 a_17685_3840.n49 10.625
R581 a_17685_3840.n49 a_17685_3840.n48 10.625
R582 a_17685_3840.n48 a_17685_3840.n47 10.625
R583 a_17685_3840.n47 a_17685_3840.n46 10.625
R584 a_17685_3840.n46 a_17685_3840.n45 10.625
R585 a_17685_3840.n45 a_17685_3840.n44 10.625
R586 a_17685_3840.n44 a_17685_3840.t19 8.716
R587 a_17685_3840.n45 a_17685_3840.t25 8.716
R588 a_17685_3840.n46 a_17685_3840.t34 8.716
R589 a_17685_3840.n47 a_17685_3840.t40 8.716
R590 a_17685_3840.n48 a_17685_3840.t17 8.716
R591 a_17685_3840.n49 a_17685_3840.t23 8.716
R592 a_17685_3840.n50 a_17685_3840.t32 8.716
R593 a_17685_3840.n51 a_17685_3840.t30 8.716
R594 a_17685_3840.n52 a_17685_3840.t37 8.716
R595 a_17685_3840.n53 a_17685_3840.t45 8.716
R596 a_17685_3840.n2 a_17685_3840.t51 8.713
R597 a_17685_3840.n3 a_17685_3840.t56 8.713
R598 a_17685_3840.n4 a_17685_3840.t64 8.713
R599 a_17685_3840.n5 a_17685_3840.t20 8.713
R600 a_17685_3840.n6 a_17685_3840.t48 8.713
R601 a_17685_3840.n7 a_17685_3840.t53 8.713
R602 a_17685_3840.n8 a_17685_3840.t60 8.713
R603 a_17685_3840.n9 a_17685_3840.t58 8.713
R604 a_17685_3840.n10 a_17685_3840.t63 8.713
R605 a_17685_3840.n11 a_17685_3840.t22 8.713
R606 a_17685_3840.n13 a_17685_3840.t42 8.708
R607 a_17685_3840.n14 a_17685_3840.t49 8.708
R608 a_17685_3840.n15 a_17685_3840.t55 8.708
R609 a_17685_3840.n16 a_17685_3840.t61 8.708
R610 a_17685_3840.n17 a_17685_3840.t18 8.708
R611 a_17685_3840.n18 a_17685_3840.t24 8.708
R612 a_17685_3840.n19 a_17685_3840.t33 8.708
R613 a_17685_3840.n20 a_17685_3840.t31 8.708
R614 a_17685_3840.n21 a_17685_3840.t38 8.708
R615 a_17685_3840.n22 a_17685_3840.t46 8.708
R616 a_17685_3840.n42 a_17685_3840.t52 8.704
R617 a_17685_3840.n33 a_17685_3840.t57 8.704
R618 a_17685_3840.n34 a_17685_3840.t62 8.704
R619 a_17685_3840.n35 a_17685_3840.t21 8.704
R620 a_17685_3840.n36 a_17685_3840.t28 8.704
R621 a_17685_3840.n37 a_17685_3840.t29 8.704
R622 a_17685_3840.n38 a_17685_3840.t36 8.704
R623 a_17685_3840.n39 a_17685_3840.t44 8.704
R624 a_17685_3840.n40 a_17685_3840.t41 8.704
R625 a_17685_3840.n41 a_17685_3840.t47 8.704
R626 a_17685_3840.n23 a_17685_3840.n22 8.14
R627 a_17685_3840.n43 a_17685_3840.n42 8.128
R628 a_17685_3840.n54 a_17685_3840.n53 8.116
R629 a_17685_3840.n12 a_17685_3840.n11 8.112
R630 a_14266_8900.t16 a_14266_8900.t25 1273.78
R631 a_14266_8900.n3 a_14266_8900.t54 193.916
R632 a_14266_8900.t54 a_14266_8900.t21 113.753
R633 a_14266_8900.t54 a_14266_8900.t11 113.753
R634 a_14266_8900.t54 a_14266_8900.t32 113.753
R635 a_14266_8900.t54 a_14266_8900.t41 113.753
R636 a_14266_8900.t54 a_14266_8900.t52 113.753
R637 a_14266_8900.t54 a_14266_8900.t50 113.753
R638 a_14266_8900.t54 a_14266_8900.t59 113.753
R639 a_14266_8900.t54 a_14266_8900.t18 113.753
R640 a_14266_8900.n2 a_14266_8900.t8 113.753
R641 a_14266_8900.n2 a_14266_8900.t48 113.753
R642 a_14266_8900.n2 a_14266_8900.t42 113.753
R643 a_14266_8900.n2 a_14266_8900.t55 113.753
R644 a_14266_8900.n0 a_14266_8900.t17 113.753
R645 a_14266_8900.n0 a_14266_8900.t34 113.753
R646 a_14266_8900.n1 a_14266_8900.t45 113.753
R647 a_14266_8900.n1 a_14266_8900.t39 113.753
R648 a_14266_8900.n1 a_14266_8900.t13 113.753
R649 a_14266_8900.n1 a_14266_8900.t5 113.753
R650 a_14266_8900.n1 a_14266_8900.t29 113.753
R651 a_14266_8900.n0 a_14266_8900.t23 113.753
R652 a_14266_8900.n0 a_14266_8900.t53 113.753
R653 a_14266_8900.n0 a_14266_8900.t51 113.753
R654 a_14266_8900.n0 a_14266_8900.t60 113.753
R655 a_14266_8900.t47 a_14266_8900.t20 113.753
R656 a_14266_8900.t47 a_14266_8900.t9 113.753
R657 a_14266_8900.t47 a_14266_8900.t49 113.753
R658 a_14266_8900.t47 a_14266_8900.t43 113.753
R659 a_14266_8900.t47 a_14266_8900.t56 113.753
R660 a_14266_8900.n0 a_14266_8900.t19 113.753
R661 a_14266_8900.t47 a_14266_8900.t35 113.753
R662 a_14266_8900.t47 a_14266_8900.t46 113.753
R663 a_14266_8900.t47 a_14266_8900.t40 113.753
R664 a_14266_8900.t47 a_14266_8900.t14 113.753
R665 a_14266_8900.t47 a_14266_8900.t6 113.753
R666 a_14266_8900.t47 a_14266_8900.t30 113.753
R667 a_14266_8900.n0 a_14266_8900.t24 113.753
R668 a_14266_8900.n0 a_14266_8900.t2 113.753
R669 a_14266_8900.n0 a_14266_8900.t61 113.753
R670 a_14266_8900.t47 a_14266_8900.t27 113.753
R671 a_14266_8900.t47 a_14266_8900.t36 113.753
R672 a_14266_8900.t47 a_14266_8900.t31 113.753
R673 a_14266_8900.t47 a_14266_8900.t58 113.753
R674 a_14266_8900.t47 a_14266_8900.t57 113.753
R675 a_14266_8900.t47 a_14266_8900.t7 113.753
R676 a_14266_8900.t54 a_14266_8900.t22 113.753
R677 a_14266_8900.t54 a_14266_8900.t15 113.753
R678 a_14266_8900.t54 a_14266_8900.t33 113.753
R679 a_14266_8900.t54 a_14266_8900.t44 113.753
R680 a_14266_8900.t47 a_14266_8900.t38 113.753
R681 a_14266_8900.t47 a_14266_8900.t12 113.753
R682 a_14266_8900.t47 a_14266_8900.t4 113.753
R683 a_14266_8900.t47 a_14266_8900.t28 113.753
R684 a_14266_8900.t54 a_14266_8900.t37 113.753
R685 a_14266_8900.t54 a_14266_8900.t10 113.753
R686 a_14266_8900.t54 a_14266_8900.t3 113.753
R687 a_14266_8900.t54 a_14266_8900.t26 113.753
R688 a_14266_8900.t0 a_14266_8900.n4 57.619
R689 a_14266_8900.n4 a_14266_8900.n3 43.122
R690 a_14266_8900.n3 a_14266_8900.t1 28.571
R691 a_14266_8900.n4 a_14266_8900.t16 10.022
R692 a_14266_8900.t54 a_14266_8900.n0 5.834
R693 a_14266_8900.t47 a_14266_8900.n1 2.869
R694 a_14266_8900.t54 a_14266_8900.t47 2.813
R695 a_14266_8900.t47 a_14266_8900.n2 2.586
R696 a_52052_20860.t9 a_52052_20860.n16 2527.24
R697 a_52052_20860.n8 a_52052_20860.t17 212.622
R698 a_52052_20860.n5 a_52052_20860.t7 212.622
R699 a_52052_20860.n12 a_52052_20860.n10 208.271
R700 a_52052_20860.n2 a_52052_20860.n0 208.271
R701 a_52052_20860.n14 a_52052_20860.n12 208.271
R702 a_52052_20860.n9 a_52052_20860.n8 208.271
R703 a_52052_20860.n4 a_52052_20860.n2 208.271
R704 a_52052_20860.n6 a_52052_20860.n5 208.271
R705 a_52052_20860.n7 a_52052_20860.n6 122.265
R706 a_52052_20860.n15 a_52052_20860.n14 121.297
R707 a_52052_20860.n7 a_52052_20860.n4 63.478
R708 a_52052_20860.n15 a_52052_20860.n9 63.217
R709 a_52052_20860.n16 a_52052_20860.n7 38.746
R710 a_52052_20860.n16 a_52052_20860.n15 15.694
R711 a_52052_20860.n8 a_52052_20860.t14 4.351
R712 a_52052_20860.n9 a_52052_20860.t11 4.351
R713 a_52052_20860.n5 a_52052_20860.t4 4.351
R714 a_52052_20860.n6 a_52052_20860.t1 4.351
R715 a_52052_20860.n10 a_52052_20860.t13 4.35
R716 a_52052_20860.n10 a_52052_20860.t18 4.35
R717 a_52052_20860.n11 a_52052_20860.t10 4.35
R718 a_52052_20860.n11 a_52052_20860.t16 4.35
R719 a_52052_20860.n13 a_52052_20860.t15 4.35
R720 a_52052_20860.n13 a_52052_20860.t12 4.35
R721 a_52052_20860.n0 a_52052_20860.t3 4.35
R722 a_52052_20860.n0 a_52052_20860.t8 4.35
R723 a_52052_20860.n1 a_52052_20860.t0 4.35
R724 a_52052_20860.n1 a_52052_20860.t6 4.35
R725 a_52052_20860.n3 a_52052_20860.t5 4.35
R726 a_52052_20860.n3 a_52052_20860.t2 4.35
R727 a_52052_20860.n14 a_52052_20860.n13 0.001
R728 a_52052_20860.n12 a_52052_20860.n11 0.001
R729 a_52052_20860.n4 a_52052_20860.n3 0.001
R730 a_52052_20860.n2 a_52052_20860.n1 0.001
R731 a_56334_20860.n0 a_56334_20860.t2 171.564
R732 a_56334_20860.n0 a_56334_20860.t1 171.563
R733 a_56334_20860.t0 a_56334_20860.n0 171.52
R734 a_23156_5032.n0 a_23156_5032.t7 365.308
R735 a_23156_5032.n4 a_23156_5032.t2 93.107
R736 a_23156_5032.n5 a_23156_5032.n4 75.71
R737 a_23156_5032.n3 a_23156_5032.n2 75.707
R738 a_23156_5032.n2 a_23156_5032.n1 75.707
R739 a_23156_5032.n1 a_23156_5032.n0 75.707
R740 a_23156_5032.n5 a_23156_5032.n3 75.706
R741 a_23156_5032.t6 a_23156_5032.n5 17.401
R742 a_23156_5032.n0 a_23156_5032.t3 17.401
R743 a_23156_5032.n1 a_23156_5032.t0 17.401
R744 a_23156_5032.n2 a_23156_5032.t5 17.401
R745 a_23156_5032.n3 a_23156_5032.t1 17.401
R746 a_23156_5032.n4 a_23156_5032.t4 17.401
R747 a_23436_16644.t46 a_23436_16644.t43 1273.78
R748 a_23436_16644.n3 a_23436_16644.t0 1158.7
R749 a_23436_16644.n3 a_23436_16644.t60 169.095
R750 a_23436_16644.t60 a_23436_16644.t45 113.753
R751 a_23436_16644.t60 a_23436_16644.t5 113.753
R752 a_23436_16644.t60 a_23436_16644.t21 113.753
R753 a_23436_16644.t60 a_23436_16644.t20 113.753
R754 a_23436_16644.t60 a_23436_16644.t2 113.753
R755 a_23436_16644.t60 a_23436_16644.t17 113.753
R756 a_23436_16644.t60 a_23436_16644.t37 113.753
R757 a_23436_16644.t60 a_23436_16644.t33 113.753
R758 a_23436_16644.n2 a_23436_16644.t44 113.753
R759 a_23436_16644.n2 a_23436_16644.t59 113.753
R760 a_23436_16644.n2 a_23436_16644.t14 113.753
R761 a_23436_16644.n2 a_23436_16644.t32 113.753
R762 a_23436_16644.n0 a_23436_16644.t10 113.753
R763 a_23436_16644.n0 a_23436_16644.t28 113.753
R764 a_23436_16644.n1 a_23436_16644.t26 113.753
R765 a_23436_16644.n1 a_23436_16644.t34 113.753
R766 a_23436_16644.n1 a_23436_16644.t47 113.753
R767 a_23436_16644.n1 a_23436_16644.t6 113.753
R768 a_23436_16644.n1 a_23436_16644.t24 113.753
R769 a_23436_16644.n0 a_23436_16644.t50 113.753
R770 a_23436_16644.n0 a_23436_16644.t22 113.753
R771 a_23436_16644.n0 a_23436_16644.t40 113.753
R772 a_23436_16644.n0 a_23436_16644.t58 113.753
R773 a_23436_16644.t12 a_23436_16644.t56 113.753
R774 a_23436_16644.t12 a_23436_16644.t8 113.753
R775 a_23436_16644.t12 a_23436_16644.t18 113.753
R776 a_23436_16644.t12 a_23436_16644.t38 113.753
R777 a_23436_16644.t12 a_23436_16644.t54 113.753
R778 a_23436_16644.n0 a_23436_16644.t11 113.753
R779 a_23436_16644.t12 a_23436_16644.t29 113.753
R780 a_23436_16644.t12 a_23436_16644.t27 113.753
R781 a_23436_16644.t12 a_23436_16644.t35 113.753
R782 a_23436_16644.t12 a_23436_16644.t48 113.753
R783 a_23436_16644.t12 a_23436_16644.t7 113.753
R784 a_23436_16644.t12 a_23436_16644.t25 113.753
R785 a_23436_16644.n0 a_23436_16644.t51 113.753
R786 a_23436_16644.n0 a_23436_16644.t23 113.753
R787 a_23436_16644.n0 a_23436_16644.t41 113.753
R788 a_23436_16644.t12 a_23436_16644.t61 113.753
R789 a_23436_16644.t12 a_23436_16644.t57 113.753
R790 a_23436_16644.t12 a_23436_16644.t9 113.753
R791 a_23436_16644.t12 a_23436_16644.t19 113.753
R792 a_23436_16644.t12 a_23436_16644.t39 113.753
R793 a_23436_16644.t12 a_23436_16644.t55 113.753
R794 a_23436_16644.t60 a_23436_16644.t15 113.753
R795 a_23436_16644.t60 a_23436_16644.t36 113.753
R796 a_23436_16644.t60 a_23436_16644.t53 113.753
R797 a_23436_16644.t60 a_23436_16644.t52 113.753
R798 a_23436_16644.t12 a_23436_16644.t4 113.753
R799 a_23436_16644.t12 a_23436_16644.t13 113.753
R800 a_23436_16644.t12 a_23436_16644.t31 113.753
R801 a_23436_16644.t12 a_23436_16644.t49 113.753
R802 a_23436_16644.t60 a_23436_16644.t30 113.753
R803 a_23436_16644.t60 a_23436_16644.t42 113.753
R804 a_23436_16644.t60 a_23436_16644.t3 113.753
R805 a_23436_16644.t60 a_23436_16644.t16 113.753
R806 a_23436_16644.t1 a_23436_16644.n3 59.624
R807 a_23436_16644.t60 a_23436_16644.t46 6.578
R808 a_23436_16644.t60 a_23436_16644.n0 5.834
R809 a_23436_16644.t12 a_23436_16644.n1 2.869
R810 a_23436_16644.t12 a_23436_16644.n2 2.586
R811 a_23436_16644.t60 a_23436_16644.t12 2.576
R812 a_25778_4988.n0 a_25778_4988.t7 334.707
R813 a_25778_4988.n4 a_25778_4988.t2 93.107
R814 a_25778_4988.n5 a_25778_4988.n4 75.71
R815 a_25778_4988.n3 a_25778_4988.n2 75.707
R816 a_25778_4988.n2 a_25778_4988.n1 75.707
R817 a_25778_4988.n1 a_25778_4988.n0 75.707
R818 a_25778_4988.n5 a_25778_4988.n3 75.706
R819 a_25778_4988.t6 a_25778_4988.n5 17.401
R820 a_25778_4988.n0 a_25778_4988.t3 17.401
R821 a_25778_4988.n1 a_25778_4988.t0 17.401
R822 a_25778_4988.n2 a_25778_4988.t5 17.401
R823 a_25778_4988.n3 a_25778_4988.t1 17.401
R824 a_25778_4988.n4 a_25778_4988.t4 17.401
R825 Fvco.t28 Fvco.t8 1273.78
R826 Fvco.t28 Fvco.n3 132.569
R827 Fvco.t4 Fvco.t25 113.753
R828 Fvco.t4 Fvco.t24 113.753
R829 Fvco.t4 Fvco.t35 113.753
R830 Fvco.t4 Fvco.t48 113.753
R831 Fvco.n2 Fvco.t47 113.753
R832 Fvco.n2 Fvco.t23 113.753
R833 Fvco.n2 Fvco.t20 113.753
R834 Fvco.n2 Fvco.t30 113.753
R835 Fvco.n0 Fvco.t13 113.753
R836 Fvco.n0 Fvco.t27 113.753
R837 Fvco.t26 Fvco.t38 113.753
R838 Fvco.t26 Fvco.t32 113.753
R839 Fvco.t26 Fvco.t11 113.753
R840 Fvco.t26 Fvco.t6 113.753
R841 Fvco.t26 Fvco.t21 113.753
R842 Fvco.n0 Fvco.t17 113.753
R843 Fvco.n0 Fvco.t44 113.753
R844 Fvco.n0 Fvco.t42 113.753
R845 Fvco.n0 Fvco.t2 113.753
R846 Fvco.t26 Fvco.t15 113.753
R847 Fvco.t26 Fvco.t9 113.753
R848 Fvco.t26 Fvco.t40 113.753
R849 Fvco.t26 Fvco.t36 113.753
R850 Fvco.t26 Fvco.t49 113.753
R851 Fvco.n0 Fvco.t14 113.753
R852 Fvco.t26 Fvco.t29 113.753
R853 Fvco.t26 Fvco.t39 113.753
R854 Fvco.t26 Fvco.t33 113.753
R855 Fvco.t26 Fvco.t12 113.753
R856 Fvco.t26 Fvco.t7 113.753
R857 Fvco.t26 Fvco.t22 113.753
R858 Fvco.n0 Fvco.t18 113.753
R859 Fvco.n0 Fvco.t45 113.753
R860 Fvco.n0 Fvco.t43 113.753
R861 Fvco.n1 Fvco.t3 113.753
R862 Fvco.n1 Fvco.t16 113.753
R863 Fvco.n1 Fvco.t10 113.753
R864 Fvco.n1 Fvco.t41 113.753
R865 Fvco.t26 Fvco.t37 113.753
R866 Fvco.t26 Fvco.t50 113.753
R867 Fvco.t4 Fvco.t5 113.753
R868 Fvco.t4 Fvco.t34 113.753
R869 Fvco.t4 Fvco.t31 113.753
R870 Fvco.t4 Fvco.t46 113.753
R871 Fvco.t4 Fvco.t19 113.753
R872 Fvco.n3 Fvco.t0 77.367
R873 Fvco.n3 Fvco.t1 28.578
R874 Fvco.t28 Fvco.t4 5.352
R875 Fvco.t4 Fvco.t26 4.314
R876 Fvco.t4 Fvco.n0 3.605
R877 Fvco.t26 Fvco.n1 2.943
R878 Fvco.t4 Fvco.n2 2.578
R879 vbiasob.n2 vbiasob.t1 67.964
R880 vbiasob.n0 vbiasob.t3 61.399
R881 vbiasob.n0 vbiasob.t4 60.299
R882 vbiasob.n1 vbiasob.t0 18.573
R883 vbiasob.n3 vbiasob.n2 12.525
R884 vbiasob.n1 vbiasob.t2 5.717
R885 vbiasob.n2 vbiasob.n1 1.012
R886 vbiasob.n3 vbiasob.n0 0.614
R887 vbiasob vbiasob.n3 0.484
R888 a_56272_15934.t1 a_56272_15934.t0 409.924
R889 vbiasbuffer.n0 vbiasbuffer.t1 136.915
R890 vbiasbuffer.n1 vbiasbuffer.t4 125.304
R891 vbiasbuffer.n1 vbiasbuffer.t3 120.586
R892 vbiasbuffer.n0 vbiasbuffer.t0 22.405
R893 vbiasbuffer vbiasbuffer.n0 15.01
R894 vbiasbuffer.n0 vbiasbuffer.t2 5.719
R895 vbiasbuffer vbiasbuffer.n1 0.631
R896 a_57726_5786.n0 a_57726_5786.t2 85.561
R897 a_57726_5786.n1 a_57726_5786.t0 85.561
R898 a_57726_5786.n0 a_57726_5786.t5 39.685
R899 a_57726_5786.n1 a_57726_5786.t4 17.517
R900 a_57726_5786.t3 a_57726_5786.n3 5.8
R901 a_57726_5786.n3 a_57726_5786.t1 5.8
R902 a_57726_5786.n3 a_57726_5786.n2 0.736
R903 a_57726_5786.n2 a_57726_5786.n0 0.231
R904 a_57726_5786.n2 a_57726_5786.n1 0.206
R905 a_28578_5014.n5 a_28578_5014.t7 265.844
R906 a_28578_5014.n0 a_28578_5014.t5 93.107
R907 a_28578_5014.n5 a_28578_5014.n4 75.71
R908 a_28578_5014.n1 a_28578_5014.n0 75.707
R909 a_28578_5014.n2 a_28578_5014.n1 75.707
R910 a_28578_5014.n3 a_28578_5014.n2 75.707
R911 a_28578_5014.n4 a_28578_5014.n3 75.707
R912 a_28578_5014.t6 a_28578_5014.n5 17.401
R913 a_28578_5014.n4 a_28578_5014.t3 17.401
R914 a_28578_5014.n3 a_28578_5014.t1 17.401
R915 a_28578_5014.n2 a_28578_5014.t4 17.401
R916 a_28578_5014.n1 a_28578_5014.t2 17.401
R917 a_28578_5014.n0 a_28578_5014.t0 17.401
R918 a_50583_13108.n0 a_50583_13108.t2 1776.66
R919 a_50583_13108.n0 a_50583_13108.t1 171.607
R920 a_50583_13108.t0 a_50583_13108.n0 171.607
R921 vinit.n9 vinit.t44 56.95
R922 vinit.n11 vinit.t42 56.876
R923 vinit.n12 vinit.t43 56.876
R924 vinit.n10 vinit.t40 56.876
R925 vinit.n9 vinit.t41 56.876
R926 vinit.n15 vinit.n14 32.801
R927 vinit.n15 vinit.t37 7.425
R928 vinit.n34 vinit.t24 7.425
R929 vinit.n32 vinit.t32 5.713
R930 vinit.n32 vinit.t30 5.713
R931 vinit.n30 vinit.t36 5.713
R932 vinit.n30 vinit.t21 5.713
R933 vinit.n28 vinit.t23 5.713
R934 vinit.n28 vinit.t29 5.713
R935 vinit.n26 vinit.t28 5.713
R936 vinit.n26 vinit.t35 5.713
R937 vinit.n24 vinit.t38 5.713
R938 vinit.n24 vinit.t22 5.713
R939 vinit.n22 vinit.t27 5.713
R940 vinit.n22 vinit.t26 5.713
R941 vinit.n20 vinit.t33 5.713
R942 vinit.n20 vinit.t31 5.713
R943 vinit.n18 vinit.t20 5.713
R944 vinit.n18 vinit.t25 5.713
R945 vinit.n16 vinit.t34 5.713
R946 vinit.n16 vinit.t39 5.713
R947 vinit.n45 vinit.t3 5.244
R948 vinit.n35 vinit.t16 5.244
R949 vinit.n0 vinit.t1 3.48
R950 vinit.n0 vinit.t8 3.48
R951 vinit.n1 vinit.t7 3.48
R952 vinit.n1 vinit.t14 3.48
R953 vinit.n2 vinit.t0 3.48
R954 vinit.n2 vinit.t19 3.48
R955 vinit.n3 vinit.t6 3.48
R956 vinit.n3 vinit.t5 3.48
R957 vinit.n4 vinit.t12 3.48
R958 vinit.n4 vinit.t15 3.48
R959 vinit.n5 vinit.t18 3.48
R960 vinit.n5 vinit.t4 3.48
R961 vinit.n6 vinit.t2 3.48
R962 vinit.n6 vinit.t9 3.48
R963 vinit.n7 vinit.t13 3.48
R964 vinit.n7 vinit.t17 3.48
R965 vinit.n8 vinit.t11 3.48
R966 vinit.n8 vinit.t10 3.48
R967 vinit.n41 vinit.n3 1.766
R968 vinit.n44 vinit.n0 1.766
R969 vinit.n38 vinit.n6 1.766
R970 vinit.n37 vinit.n7 1.764
R971 vinit.n40 vinit.n4 1.762
R972 vinit.n42 vinit.n2 1.761
R973 vinit.n39 vinit.n5 1.758
R974 vinit.n43 vinit.n1 1.758
R975 vinit.n36 vinit.n8 1.754
R976 vinit.n23 vinit.n22 1.714
R977 vinit.n17 vinit.n16 1.714
R978 vinit.n29 vinit.n28 1.714
R979 vinit.n31 vinit.n30 1.712
R980 vinit.n25 vinit.n24 1.71
R981 vinit.n21 vinit.n20 1.709
R982 vinit.n27 vinit.n26 1.706
R983 vinit.n19 vinit.n18 1.706
R984 vinit.n33 vinit.n32 1.702
R985 vinit.n14 vinit.n13 0.322
R986 vinit.n35 vinit.n34 0.295
R987 vinit vinit.n45 0.112
R988 vinit.n12 vinit.n11 0.073
R989 vinit.n10 vinit.n9 0.073
R990 vinit.n13 vinit.n12 0.051
R991 vinit.n34 vinit.n33 0.032
R992 vinit.n40 vinit.n39 0.031
R993 vinit.n27 vinit.n25 0.031
R994 vinit.n43 vinit.n42 0.031
R995 vinit.n21 vinit.n19 0.031
R996 vinit.n37 vinit.n36 0.031
R997 vinit.n33 vinit.n31 0.031
R998 vinit.n36 vinit.n35 0.031
R999 vinit.n44 vinit.n43 0.03
R1000 vinit.n19 vinit.n17 0.03
R1001 vinit.n45 vinit.n44 0.03
R1002 vinit.n17 vinit.n15 0.03
R1003 vinit.n38 vinit.n37 0.03
R1004 vinit.n31 vinit.n29 0.03
R1005 vinit.n41 vinit.n40 0.03
R1006 vinit.n25 vinit.n23 0.03
R1007 vinit.n42 vinit.n41 0.03
R1008 vinit.n23 vinit.n21 0.03
R1009 vinit.n39 vinit.n38 0.03
R1010 vinit.n29 vinit.n27 0.03
R1011 vinit.n13 vinit.n10 0.022
R1012 a_27762_11446.t11 a_27762_11446.t48 1273.78
R1013 a_27762_11446.t47 a_27762_11446.t13 113.753
R1014 a_27762_11446.t47 a_27762_11446.t23 113.753
R1015 a_27762_11446.t47 a_27762_11446.t39 113.753
R1016 a_27762_11446.t47 a_27762_11446.t56 113.753
R1017 a_27762_11446.t47 a_27762_11446.t45 113.753
R1018 a_27762_11446.t47 a_27762_11446.t60 113.753
R1019 a_27762_11446.t47 a_27762_11446.t9 113.753
R1020 a_27762_11446.t47 a_27762_11446.t30 113.753
R1021 a_27762_11446.n2 a_27762_11446.t25 113.753
R1022 a_27762_11446.n2 a_27762_11446.t37 113.753
R1023 a_27762_11446.n2 a_27762_11446.t53 113.753
R1024 a_27762_11446.n2 a_27762_11446.t7 113.753
R1025 a_27762_11446.n0 a_27762_11446.t28 113.753
R1026 a_27762_11446.n0 a_27762_11446.t41 113.753
R1027 a_27762_11446.n1 a_27762_11446.t58 113.753
R1028 a_27762_11446.n1 a_27762_11446.t51 113.753
R1029 a_27762_11446.n1 a_27762_11446.t5 113.753
R1030 a_27762_11446.n1 a_27762_11446.t20 113.753
R1031 a_27762_11446.n1 a_27762_11446.t35 113.753
R1032 a_27762_11446.n0 a_27762_11446.t15 113.753
R1033 a_27762_11446.n0 a_27762_11446.t46 113.753
R1034 a_27762_11446.n0 a_27762_11446.t61 113.753
R1035 a_27762_11446.n0 a_27762_11446.t10 113.753
R1036 a_27762_11446.t21 a_27762_11446.t31 113.753
R1037 a_27762_11446.t21 a_27762_11446.t26 113.753
R1038 a_27762_11446.t21 a_27762_11446.t38 113.753
R1039 a_27762_11446.t21 a_27762_11446.t54 113.753
R1040 a_27762_11446.t21 a_27762_11446.t8 113.753
R1041 a_27762_11446.n0 a_27762_11446.t29 113.753
R1042 a_27762_11446.t21 a_27762_11446.t42 113.753
R1043 a_27762_11446.t21 a_27762_11446.t59 113.753
R1044 a_27762_11446.t21 a_27762_11446.t52 113.753
R1045 a_27762_11446.t21 a_27762_11446.t6 113.753
R1046 a_27762_11446.t21 a_27762_11446.t22 113.753
R1047 a_27762_11446.t21 a_27762_11446.t36 113.753
R1048 a_27762_11446.n0 a_27762_11446.t16 113.753
R1049 a_27762_11446.n0 a_27762_11446.t3 113.753
R1050 a_27762_11446.n0 a_27762_11446.t17 113.753
R1051 a_27762_11446.t21 a_27762_11446.t32 113.753
R1052 a_27762_11446.t21 a_27762_11446.t44 113.753
R1053 a_27762_11446.t21 a_27762_11446.t43 113.753
R1054 a_27762_11446.t21 a_27762_11446.t55 113.753
R1055 a_27762_11446.t21 a_27762_11446.t12 113.753
R1056 a_27762_11446.t21 a_27762_11446.t24 113.753
R1057 a_27762_11446.t47 a_27762_11446.t14 113.753
R1058 a_27762_11446.t47 a_27762_11446.t27 113.753
R1059 a_27762_11446.t47 a_27762_11446.t40 113.753
R1060 a_27762_11446.t47 a_27762_11446.t57 113.753
R1061 a_27762_11446.t21 a_27762_11446.t50 113.753
R1062 a_27762_11446.t21 a_27762_11446.t4 113.753
R1063 a_27762_11446.t21 a_27762_11446.t19 113.753
R1064 a_27762_11446.t21 a_27762_11446.t34 113.753
R1065 a_27762_11446.t47 a_27762_11446.t49 113.753
R1066 a_27762_11446.t47 a_27762_11446.t2 113.753
R1067 a_27762_11446.t47 a_27762_11446.t18 113.753
R1068 a_27762_11446.t47 a_27762_11446.t33 113.753
R1069 a_27762_11446.n4 a_27762_11446.n3 88.886
R1070 a_27762_11446.n4 a_27762_11446.t0 81.996
R1071 a_27762_11446.t1 a_27762_11446.n4 59.267
R1072 a_27762_11446.t47 a_27762_11446.n0 5.834
R1073 a_27762_11446.n3 a_27762_11446.t11 4.994
R1074 a_27762_11446.n3 a_27762_11446.t47 4.809
R1075 a_27762_11446.t21 a_27762_11446.n1 2.869
R1076 a_27762_11446.t47 a_27762_11446.t21 2.8
R1077 a_27762_11446.t21 a_27762_11446.n2 2.586
R1078 a_49932_4124.t1 a_49932_4124.t2 33.597
R1079 a_49932_4124.t0 a_49932_4124.t1 13.614
R1080 a_49932_4124.t1 a_49932_4124.t3 11.692
R1081 a_44752_16348.t4 a_44752_16348.n2 349.137
R1082 a_44752_16348.n1 a_44752_16348.t1 197.553
R1083 a_44752_16348.n0 a_44752_16348.t2 178.539
R1084 a_44752_16348.n0 a_44752_16348.t3 122.603
R1085 a_44752_16348.n1 a_44752_16348.t0 114.713
R1086 a_44752_16348.n2 a_44752_16348.n0 95.215
R1087 a_44752_16348.n2 a_44752_16348.n1 26.034
R1088 a_51138_19904.n0 a_51138_19904.t2 171.567
R1089 a_51138_19904.t0 a_51138_19904.n0 171.564
R1090 a_51138_19904.n0 a_51138_19904.t1 171.52
R1091 a_14832_12082.n1 a_14832_12082.t3 434.515
R1092 a_14832_12082.n0 a_14832_12082.t2 217.163
R1093 a_14832_12082.t1 a_14832_12082.n1 52.152
R1094 a_14832_12082.n0 a_14832_12082.t0 3.106
R1095 a_14832_12082.n1 a_14832_12082.n0 0.908
R1096 CLK_BY_4_IPH_BAR.n3 CLK_BY_4_IPH_BAR.t8 449.587
R1097 CLK_BY_4_IPH_BAR.n3 CLK_BY_4_IPH_BAR.t3 402.739
R1098 CLK_BY_4_IPH_BAR.n7 CLK_BY_4_IPH_BAR.t6 333.651
R1099 CLK_BY_4_IPH_BAR.n7 CLK_BY_4_IPH_BAR.t7 297.233
R1100 CLK_BY_4_IPH_BAR.n2 CLK_BY_4_IPH_BAR.t4 270.989
R1101 CLK_BY_4_IPH_BAR.n2 CLK_BY_4_IPH_BAR.t5 227.612
R1102 CLK_BY_4_IPH_BAR.n4 CLK_BY_4_IPH_BAR.n2 199.119
R1103 CLK_BY_4_IPH_BAR.n5 CLK_BY_4_IPH_BAR.n4 138.541
R1104 CLK_BY_4_IPH_BAR.n5 CLK_BY_4_IPH_BAR.t2 98.31
R1105 CLK_BY_4_IPH_BAR.n0 CLK_BY_4_IPH_BAR.t1 92.047
R1106 CLK_BY_4_IPH_BAR.n8 CLK_BY_4_IPH_BAR.n7 70.234
R1107 CLK_BY_4_IPH_BAR.n0 CLK_BY_4_IPH_BAR.t0 61.427
R1108 CLK_BY_4_IPH_BAR.n4 CLK_BY_4_IPH_BAR.n3 38.57
R1109 CLK_BY_4_IPH_BAR.n6 CLK_BY_4_IPH_BAR.n5 1.254
R1110 CLK_BY_4_IPH_BAR.n6 CLK_BY_4_IPH_BAR.n1 0.057
R1111 CLK_BY_4_IPH_BAR.n1 CLK_BY_4_IPH_BAR.n0 0.055
R1112 CLK_BY_4_IPH_BAR CLK_BY_4_IPH_BAR.n8 0.016
R1113 CLK_BY_4_IPH_BAR CLK_BY_4_IPH_BAR.n6 0.012
R1114 a_23160_10936.n5 a_23160_10936.t7 391.966
R1115 a_23160_10936.n0 a_23160_10936.t5 93.107
R1116 a_23160_10936.n5 a_23160_10936.n4 75.709
R1117 a_23160_10936.n1 a_23160_10936.n0 75.707
R1118 a_23160_10936.n2 a_23160_10936.n1 75.707
R1119 a_23160_10936.n3 a_23160_10936.n2 75.707
R1120 a_23160_10936.n4 a_23160_10936.n3 75.707
R1121 a_23160_10936.t6 a_23160_10936.n5 17.401
R1122 a_23160_10936.n4 a_23160_10936.t2 17.401
R1123 a_23160_10936.n3 a_23160_10936.t0 17.401
R1124 a_23160_10936.n2 a_23160_10936.t3 17.401
R1125 a_23160_10936.n1 a_23160_10936.t1 17.401
R1126 a_23160_10936.n0 a_23160_10936.t4 17.401
R1127 a_28438_10874.n0 a_28438_10874.t7 338.927
R1128 a_28438_10874.n4 a_28438_10874.t3 93.107
R1129 a_28438_10874.n5 a_28438_10874.n4 75.71
R1130 a_28438_10874.n1 a_28438_10874.n0 75.708
R1131 a_28438_10874.n3 a_28438_10874.n2 75.707
R1132 a_28438_10874.n2 a_28438_10874.n1 75.707
R1133 a_28438_10874.n5 a_28438_10874.n3 75.706
R1134 a_28438_10874.t6 a_28438_10874.n5 17.401
R1135 a_28438_10874.n0 a_28438_10874.t4 17.401
R1136 a_28438_10874.n1 a_28438_10874.t0 17.401
R1137 a_28438_10874.n2 a_28438_10874.t5 17.401
R1138 a_28438_10874.n3 a_28438_10874.t1 17.401
R1139 a_28438_10874.n4 a_28438_10874.t2 17.401
R1140 a_14910_6932.n1 a_14910_6932.t3 434.494
R1141 a_14910_6932.n0 a_14910_6932.t2 217.163
R1142 a_14910_6932.t1 a_14910_6932.n1 52.318
R1143 a_14910_6932.n0 a_14910_6932.t0 3.106
R1144 a_14910_6932.n1 a_14910_6932.n0 0.906
R1145 CLK_BY_2_BAR.n0 CLK_BY_2_BAR.t6 333.651
R1146 CLK_BY_2_BAR.n0 CLK_BY_2_BAR.t9 297.233
R1147 CLK_BY_2_BAR.n3 CLK_BY_2_BAR.t3 294.554
R1148 CLK_BY_2_BAR.n1 CLK_BY_2_BAR.t5 212.079
R1149 CLK_BY_2_BAR.n2 CLK_BY_2_BAR.t2 212.079
R1150 CLK_BY_2_BAR.n3 CLK_BY_2_BAR.t4 211.008
R1151 CLK_BY_2_BAR.n1 CLK_BY_2_BAR.t8 139.779
R1152 CLK_BY_2_BAR.n2 CLK_BY_2_BAR.t7 139.779
R1153 CLK_BY_2_BAR.n4 CLK_BY_2_BAR.t1 102.408
R1154 CLK_BY_2_BAR.n6 CLK_BY_2_BAR.n2 68.902
R1155 CLK_BY_2_BAR.n2 CLK_BY_2_BAR.n1 61.345
R1156 CLK_BY_2_BAR.n5 CLK_BY_2_BAR.t0 54.537
R1157 CLK_BY_2_BAR CLK_BY_2_BAR.n0 49.8
R1158 CLK_BY_2_BAR CLK_BY_2_BAR.n6 19.824
R1159 CLK_BY_2_BAR.n4 CLK_BY_2_BAR.n3 12.821
R1160 CLK_BY_2_BAR.n5 CLK_BY_2_BAR.n4 3.763
R1161 CLK_BY_2_BAR.n6 CLK_BY_2_BAR.n5 0.621
R1162 a_26016_10878.n0 a_26016_10878.t0 305.609
R1163 a_26016_10878.t6 a_26016_10878.n5 93.107
R1164 a_26016_10878.n1 a_26016_10878.n0 75.708
R1165 a_26016_10878.n5 a_26016_10878.n4 75.707
R1166 a_26016_10878.n4 a_26016_10878.n3 75.707
R1167 a_26016_10878.n3 a_26016_10878.n2 75.707
R1168 a_26016_10878.n2 a_26016_10878.n1 75.707
R1169 a_26016_10878.n0 a_26016_10878.t7 17.401
R1170 a_26016_10878.n1 a_26016_10878.t3 17.401
R1171 a_26016_10878.n2 a_26016_10878.t1 17.401
R1172 a_26016_10878.n3 a_26016_10878.t4 17.401
R1173 a_26016_10878.n4 a_26016_10878.t2 17.401
R1174 a_26016_10878.n5 a_26016_10878.t5 17.401
R1175 a_77280_24640.n1 a_77280_24640.t3 263.373
R1176 a_77280_24640.t0 a_77280_24640.n2 61.061
R1177 a_77280_24640.n0 a_77280_24640.t4 14.065
R1178 a_77280_24640.n0 a_77280_24640.t2 4.819
R1179 a_77280_24640.n2 a_77280_24640.n0 2.726
R1180 a_77280_24640.n1 a_77280_24640.t1 1.368
R1181 a_77280_24640.n2 a_77280_24640.n1 0.571
R1182 a_77254_23336.t6 a_77254_23336.n3 95.488
R1183 a_77254_23336.n0 a_77254_23336.t3 52.208
R1184 a_77254_23336.n3 a_77254_23336.n2 13.658
R1185 a_77254_23336.n3 a_77254_23336.t0 4.572
R1186 a_77254_23336.n1 a_77254_23336.t2 3.848
R1187 a_77254_23336.n0 a_77254_23336.t5 1.482
R1188 a_77254_23336.n2 a_77254_23336.n1 1.338
R1189 a_77254_23336.n1 a_77254_23336.t4 0.701
R1190 a_77254_23336.n2 a_77254_23336.n0 0.15
R1191 a_77254_23336.t0 a_77254_23336.t1 0.049
R1192 a_54448_7822.t1 a_54448_7822.t0 184.89
R1193 a_24410_25128.n1 a_24410_25128.t3 434.509
R1194 a_24410_25128.n0 a_24410_25128.t2 217.163
R1195 a_24410_25128.t1 a_24410_25128.n1 52.459
R1196 a_24410_25128.n0 a_24410_25128.t0 3.106
R1197 a_24410_25128.n1 a_24410_25128.n0 0.899
R1198 a_23308_802.n1 a_23308_802.t2 434.515
R1199 a_23308_802.n0 a_23308_802.t3 217.163
R1200 a_23308_802.t1 a_23308_802.n1 52.152
R1201 a_23308_802.n0 a_23308_802.t0 3.106
R1202 a_23308_802.n1 a_23308_802.n0 0.908
R1203 a_32948_24994.n1 a_32948_24994.t3 434.487
R1204 a_32948_24994.n0 a_32948_24994.t2 217.163
R1205 a_32948_24994.t1 a_32948_24994.n1 52.153
R1206 a_32948_24994.n0 a_32948_24994.t0 3.106
R1207 a_32948_24994.n1 a_32948_24994.n0 0.887
R1208 a_28790_25040.n1 a_28790_25040.t3 434.517
R1209 a_28790_25040.n0 a_28790_25040.t2 217.163
R1210 a_28790_25040.t1 a_28790_25040.n1 52.317
R1211 a_28790_25040.n0 a_28790_25040.t0 3.106
R1212 a_28790_25040.n1 a_28790_25040.n0 0.907
R1213 a_51532_4150.n1 a_51532_4150.t3 19.231
R1214 a_51532_4150.n0 a_51532_4150.t1 17.234
R1215 a_51532_4150.n2 a_51532_4150.t4 14.994
R1216 a_51532_4150.n0 a_51532_4150.t0 14.151
R1217 a_51532_4150.n1 a_51532_4150.t5 13.856
R1218 a_51532_4150.t2 a_51532_4150.n0 7.827
R1219 a_51532_4150.n1 a_51532_4150.n2 5.632
R1220 a_51532_4150.n2 a_51532_4150.t6 3.653
R1221 a_51532_4150.n0 a_51532_4150.n1 3.447
R1222 a_50032_16080.t1 a_50032_16080.t0 414.247
R1223 a_50511_16072.n4 a_50511_16072.n3 524.893
R1224 a_50511_16072.n4 a_50511_16072.t8 256.935
R1225 a_50511_16072.t7 a_50511_16072.n1 8.763
R1226 a_50511_16072.n2 a_50511_16072.t2 8.705
R1227 a_50511_16072.n1 a_50511_16072.t3 8.7
R1228 a_50511_16072.n1 a_50511_16072.t4 8.7
R1229 a_50511_16072.n0 a_50511_16072.t5 8.7
R1230 a_50511_16072.n0 a_50511_16072.t6 8.7
R1231 a_50511_16072.n3 a_50511_16072.t1 5.844
R1232 a_50511_16072.n3 a_50511_16072.t0 5.744
R1233 a_50511_16072.t8 a_50511_16072.t9 1.22
R1234 a_50511_16072.n1 a_50511_16072.n0 0.137
R1235 a_50511_16072.n0 a_50511_16072.n2 0.133
R1236 a_50511_16072.n0 a_50511_16072.n4 0.122
R1237 a_38070_8852.n1 a_38070_8852.t3 434.515
R1238 a_38070_8852.n0 a_38070_8852.t2 217.163
R1239 a_38070_8852.t1 a_38070_8852.n1 52.152
R1240 a_38070_8852.n0 a_38070_8852.t0 3.106
R1241 a_38070_8852.n1 a_38070_8852.n0 0.908
R1242 a_30384_802.n1 a_30384_802.t3 434.478
R1243 a_30384_802.n0 a_30384_802.t2 217.163
R1244 a_30384_802.t1 a_30384_802.n1 52.152
R1245 a_30384_802.n0 a_30384_802.t0 3.106
R1246 a_30384_802.n1 a_30384_802.n0 0.885
R1247 a_77598_24640.n1 a_77598_24640.t3 256.234
R1248 a_77598_24640.n0 a_77598_24640.t2 12.058
R1249 a_77598_24640.t0 a_77598_24640.n2 11.463
R1250 a_77598_24640.n0 a_77598_24640.t4 4.624
R1251 a_77598_24640.n1 a_77598_24640.t1 2.155
R1252 a_77598_24640.n2 a_77598_24640.n0 1.194
R1253 a_77598_24640.n2 a_77598_24640.n1 0.952
R1254 a_77572_23336.t4 a_77572_23336.n3 7.523
R1255 a_77572_23336.n0 a_77572_23336.t1 3.01
R1256 a_77572_23336.n1 a_77572_23336.t6 2.635
R1257 a_77572_23336.n2 a_77572_23336.t0 1.86
R1258 a_77572_23336.n3 a_77572_23336.n2 1.672
R1259 a_77572_23336.n3 a_77572_23336.n1 1.093
R1260 a_77572_23336.n0 a_77572_23336.t3 0.778
R1261 a_77572_23336.n2 a_77572_23336.t2 0.727
R1262 a_77572_23336.n1 a_77572_23336.n0 0.166
R1263 a_77572_23336.t6 a_77572_23336.t5 0.037
R1264 a_46856_21176.t0 a_46856_21176.t1 343.213
R1265 a_51138_21494.t1 a_51138_21494.t0 501.405
R1266 a_46856_19268.n0 a_46856_19268.t1 2113.41
R1267 a_46856_19268.n0 a_46856_19268.t2 171.607
R1268 a_46856_19268.t0 a_46856_19268.n0 171.607
R1269 a_51826_16054.t1 a_51826_16054.t0 445.429
R1270 a_22972_23306.n2 a_22972_23306.t1 172.018
R1271 a_22972_23306.t0 a_22972_23306.n2 171.695
R1272 a_22972_23306.n2 a_22972_23306.n1 73.17
R1273 a_22972_23306.n1 a_22972_23306.t4 28.576
R1274 a_22972_23306.n0 a_22972_23306.t2 28.565
R1275 a_22972_23306.n0 a_22972_23306.t3 28.565
R1276 a_22972_23306.n1 a_22972_23306.n0 3.497
R1277 a_54468_7504.t1 a_54468_7504.t0 178.373
R1278 b b.t0 6.636
R1279 a a.t0 4.086
C64 vbiasr gnd 146.96fF $ **FLOATING
C65 vbiasot gnd 17.09fF
C66 a_51334_14126# gnd 5.94fF
C67 a_50320_14126# gnd 7.42fF
C68 a_56602_11692# gnd 4.81fF
C69 a_55602_11692# gnd 5.68fF
C70 a_51276_14152# gnd 3.34fF
C71 a_51636_13108# gnd 8.30fF
C72 a_51041_13108# gnd 10.28fF
C73 a_50262_14152# gnd 3.87fF
C74 vbiasob gnd 11.11fF $ **FLOATING
C75 a_47760_15642# gnd 2.83fF
C76 vbiasbuffer gnd 15.97fF $ **FLOATING
C77 a_43010_16058# gnd 4.05fF
C78 a_42782_16060# gnd 4.44fF
C79 a_42574_15624# gnd 5.31fF
C80 a_42550_16062# gnd 4.20fF
C81 bb gnd 13.63fF
C82 aa gnd 15.44fF
C83 b gnd 18.62fF $ **FLOATING
C84 a gnd 14.75fF $ **FLOATING
C85 Vso8b gnd 20.82fF
C86 Vso7b gnd 14.60fF
C87 a_4226_11420# gnd 8.28fF
C88 a_4288_11534# gnd 5.07fF
C89 a_4226_11612# gnd 7.54fF
C90 a_4288_11726# gnd 6.25fF
C91 a_4226_11804# gnd 7.73fF
C92 Vso5b gnd 7.67fF
C93 Vso4b gnd 47.35fF
C94 Vso6b gnd 5.87fF
C95 a_4288_11918# gnd 5.18fF
C96 a_4226_11996# gnd 8.59fF
C97 a_4288_12110# gnd 6.31fF
C98 vout gnd 5.78fF
C99 a_4226_12188# gnd 6.34fF
C100 Fvco_By4_QPH_bar gnd 26.16fF $ **FLOATING
C101 Fvco_By4_QPH gnd 37.94fF $ **FLOATING
C102 RESET gnd 3.77fF $ **FLOATING
C103 CLK_BY_2_BAR gnd 2.66fF $ **FLOATING
C104 CLK_IN gnd 39.42fF
C105 Vso3b gnd 26.72fF
C106 Vso2b gnd 21.36fF
C107 Vso1b gnd 22.16fF
C108 vctrl gnd 12.61fF
C109 a_33808_31746# gnd 16.63fF
C110 CLK_BY_4_IPH gnd 35.38fF $ **FLOATING
C111 CLK_BY_4_IPH_BAR gnd 34.95fF $ **FLOATING
C112 vinit gnd 203.52fF $ **FLOATING
C113 a_34044_31208# gnd 377.15fF
C114 a_9354_33563# gnd 376.67fF
C115 Vdd gnd 6072.15fF
C116 a.t0 gnd 2.54fF
C117 b.t0 gnd 2.72fF
C118 a_54468_7504.t0 gnd 2.83fF
C119 a_22972_23306.n2 gnd 2.07fF $ **FLOATING
C120 a_46856_19268.n0 gnd 7.50fF $ **FLOATING
C121 a_51138_21494.t0 gnd 2.55fF
C122 a_51138_21494.t1 gnd 3.48fF
C123 a_77572_23336.t1 gnd 72.17fF
C124 a_77572_23336.t3 gnd 49.69fF
C125 a_77572_23336.n0 gnd 52.35fF $ **FLOATING
C126 a_77572_23336.t5 gnd 37.84fF $ **FLOATING
C127 a_77572_23336.t6 gnd 61.50fF $ **FLOATING
C128 a_77572_23336.n1 gnd 84.84fF $ **FLOATING
C129 a_77572_23336.t2 gnd 42.57fF
C130 a_77572_23336.t0 gnd 52.39fF
C131 a_77572_23336.n2 gnd 60.74fF $ **FLOATING
C132 a_77572_23336.n3 gnd 66.26fF $ **FLOATING
C133 a_77598_24640.t2 gnd 44.04fF $ **FLOATING
C134 a_77598_24640.t4 gnd 42.02fF $ **FLOATING
C135 a_77598_24640.n0 gnd 35.23fF $ **FLOATING
C136 a_77598_24640.t3 gnd 70.35fF $ **FLOATING
C137 a_77598_24640.t1 gnd 50.88fF $ **FLOATING
C138 a_77598_24640.n1 gnd 43.65fF $ **FLOATING
C139 a_77598_24640.n2 gnd 54.00fF $ **FLOATING
C140 a_30384_802.n0 gnd 3.14fF $ **FLOATING
C141 a_38070_8852.n0 gnd 3.65fF $ **FLOATING
C142 a_50511_16072.n0 gnd 2.15fF $ **FLOATING
C143 a_51532_4150.n1 gnd 3.34fF $ **FLOATING
C144 a_51532_4150.n2 gnd 3.10fF $ **FLOATING
C145 a_28790_25040.n0 gnd 3.75fF $ **FLOATING
C146 a_32948_24994.n0 gnd 3.11fF $ **FLOATING
C147 a_23308_802.n0 gnd 3.31fF $ **FLOATING
C148 a_24410_25128.n0 gnd 3.81fF $ **FLOATING
C149 a_54448_7822.t0 gnd 3.00fF
C150 a_77254_23336.t3 gnd 37.04fF
C151 a_77254_23336.t5 gnd 57.43fF
C152 a_77254_23336.n0 gnd 61.46fF $ **FLOATING
C153 a_77254_23336.t4 gnd 45.35fF
C154 a_77254_23336.t2 gnd 66.48fF
C155 a_77254_23336.n1 gnd 95.15fF $ **FLOATING
C156 a_77254_23336.n2 gnd 95.17fF $ **FLOATING
C157 a_77254_23336.t1 gnd 38.71fF
C158 a_77254_23336.t0 gnd 42.09fF
C159 a_77254_23336.n3 gnd 15.07fF $ **FLOATING
C160 a_77254_23336.t6 gnd 3.57fF
C161 a_77280_24640.t2 gnd 28.65fF $ **FLOATING
C162 a_77280_24640.t4 gnd 36.59fF $ **FLOATING
C163 a_77280_24640.n0 gnd 62.68fF $ **FLOATING
C164 a_77280_24640.t1 gnd 36.49fF $ **FLOATING
C165 a_77280_24640.t3 gnd 44.77fF $ **FLOATING
C166 a_77280_24640.n1 gnd 24.86fF $ **FLOATING
C167 a_77280_24640.n2 gnd 127.11fF $ **FLOATING
C168 a_77280_24640.t0 gnd 2.48fF
C169 a_14910_6932.n0 gnd 3.12fF $ **FLOATING
C170 CLK_BY_4_IPH_BAR.n5 gnd 37.30fF $ **FLOATING
C171 a_14832_12082.n0 gnd 3.86fF $ **FLOATING
C172 a_51138_19904.n0 gnd 2.56fF $ **FLOATING
C173 a_49932_4124.t1 gnd 4.56fF $ **FLOATING
C174 a_27762_11446.n0 gnd 4.89fF $ **FLOATING
C175 a_27762_11446.t47 gnd 9.88fF $ **FLOATING
C176 a_27762_11446.t21 gnd 9.88fF $ **FLOATING
C177 a_27762_11446.t11 gnd 7.39fF $ **FLOATING
C178 a_27762_11446.n3 gnd 12.90fF $ **FLOATING
C179 a_27762_11446.n4 gnd 4.16fF $ **FLOATING
C180 vinit.n14 gnd 15.21fF $ **FLOATING
C181 vinit.n15 gnd 222.87fF $ **FLOATING
C182 vinit.n34 gnd 2.69fF $ **FLOATING
C183 vinit.n35 gnd 2.72fF $ **FLOATING
C184 a_50583_13108.n0 gnd 8.05fF $ **FLOATING
C185 vbiasbuffer.n0 gnd 4.69fF $ **FLOATING
C186 vbiasob.n2 gnd 5.90fF $ **FLOATING
C187 vbiasob.n3 gnd 3.52fF $ **FLOATING
C188 Fvco.n0 gnd 3.53fF $ **FLOATING
C189 Fvco.t26 gnd 6.13fF $ **FLOATING
C190 Fvco.t4 gnd 14.39fF $ **FLOATING
C191 Fvco.t28 gnd 46.82fF $ **FLOATING
C192 Fvco.n3 gnd 4.66fF $ **FLOATING
C193 a_23436_16644.n0 gnd 4.67fF $ **FLOATING
C194 a_23436_16644.t60 gnd 10.21fF $ **FLOATING
C195 a_23436_16644.t12 gnd 8.90fF $ **FLOATING
C196 a_23436_16644.t46 gnd 6.39fF $ **FLOATING
C197 a_23436_16644.n3 gnd 3.27fF $ **FLOATING
C198 a_56334_20860.n0 gnd 2.57fF $ **FLOATING
C199 a_52052_20860.t9 gnd 3.50fF
C200 a_14266_8900.n0 gnd 4.92fF $ **FLOATING
C201 a_14266_8900.t54 gnd 9.27fF $ **FLOATING
C202 a_14266_8900.t47 gnd 9.98fF $ **FLOATING
C203 a_14266_8900.t16 gnd 12.27fF $ **FLOATING
C204 a_14266_8900.n4 gnd 10.34fF $ **FLOATING
C205 a_17685_3840.t22 gnd 2.78fF $ **FLOATING
C206 a_17685_3840.t63 gnd 2.78fF $ **FLOATING
C207 a_17685_3840.t58 gnd 2.78fF $ **FLOATING
C208 a_17685_3840.t60 gnd 2.78fF $ **FLOATING
C209 a_17685_3840.t53 gnd 2.78fF $ **FLOATING
C210 a_17685_3840.t48 gnd 2.78fF $ **FLOATING
C211 a_17685_3840.t20 gnd 2.78fF $ **FLOATING
C212 a_17685_3840.t64 gnd 2.78fF $ **FLOATING
C213 a_17685_3840.t56 gnd 2.78fF $ **FLOATING
C214 a_17685_3840.t51 gnd 2.78fF $ **FLOATING
C215 a_17685_3840.t43 gnd 6.42fF $ **FLOATING
C216 a_17685_3840.n2 gnd 11.33fF $ **FLOATING
C217 a_17685_3840.n3 gnd 7.38fF $ **FLOATING
C218 a_17685_3840.n4 gnd 7.38fF $ **FLOATING
C219 a_17685_3840.n5 gnd 7.38fF $ **FLOATING
C220 a_17685_3840.n6 gnd 7.38fF $ **FLOATING
C221 a_17685_3840.n7 gnd 7.38fF $ **FLOATING
C222 a_17685_3840.n8 gnd 7.38fF $ **FLOATING
C223 a_17685_3840.n9 gnd 7.38fF $ **FLOATING
C224 a_17685_3840.n10 gnd 7.38fF $ **FLOATING
C225 a_17685_3840.n11 gnd 6.23fF $ **FLOATING
C226 a_17685_3840.t54 gnd 3.73fF $ **FLOATING
C227 a_17685_3840.n12 gnd 7.64fF $ **FLOATING
C228 a_17685_3840.t46 gnd 2.78fF $ **FLOATING
C229 a_17685_3840.t38 gnd 2.78fF $ **FLOATING
C230 a_17685_3840.t31 gnd 2.78fF $ **FLOATING
C231 a_17685_3840.t33 gnd 2.78fF $ **FLOATING
C232 a_17685_3840.t24 gnd 2.78fF $ **FLOATING
C233 a_17685_3840.t18 gnd 2.78fF $ **FLOATING
C234 a_17685_3840.t61 gnd 2.78fF $ **FLOATING
C235 a_17685_3840.t55 gnd 2.78fF $ **FLOATING
C236 a_17685_3840.t49 gnd 2.78fF $ **FLOATING
C237 a_17685_3840.t42 gnd 2.78fF $ **FLOATING
C238 a_17685_3840.t35 gnd 6.42fF $ **FLOATING
C239 a_17685_3840.n13 gnd 11.30fF $ **FLOATING
C240 a_17685_3840.n14 gnd 7.37fF $ **FLOATING
C241 a_17685_3840.n15 gnd 7.37fF $ **FLOATING
C242 a_17685_3840.n16 gnd 7.37fF $ **FLOATING
C243 a_17685_3840.n17 gnd 7.37fF $ **FLOATING
C244 a_17685_3840.n18 gnd 7.37fF $ **FLOATING
C245 a_17685_3840.n19 gnd 7.37fF $ **FLOATING
C246 a_17685_3840.n20 gnd 7.37fF $ **FLOATING
C247 a_17685_3840.n21 gnd 7.37fF $ **FLOATING
C248 a_17685_3840.n22 gnd 6.23fF $ **FLOATING
C249 a_17685_3840.t27 gnd 3.73fF $ **FLOATING
C250 a_17685_3840.n23 gnd 5.59fF $ **FLOATING
C251 a_17685_3840.n24 gnd 6.35fF $ **FLOATING
C252 a_17685_3840.n25 gnd 3.20fF $ **FLOATING
C253 a_17685_3840.n28 gnd 2.53fF $ **FLOATING
C254 a_17685_3840.t47 gnd 2.78fF $ **FLOATING
C255 a_17685_3840.t41 gnd 2.78fF $ **FLOATING
C256 a_17685_3840.t44 gnd 2.78fF $ **FLOATING
C257 a_17685_3840.t36 gnd 2.78fF $ **FLOATING
C258 a_17685_3840.t29 gnd 2.78fF $ **FLOATING
C259 a_17685_3840.t28 gnd 2.78fF $ **FLOATING
C260 a_17685_3840.t21 gnd 2.78fF $ **FLOATING
C261 a_17685_3840.t62 gnd 2.78fF $ **FLOATING
C262 a_17685_3840.t57 gnd 2.78fF $ **FLOATING
C263 a_17685_3840.t50 gnd 6.42fF $ **FLOATING
C264 a_17685_3840.n33 gnd 11.29fF $ **FLOATING
C265 a_17685_3840.n34 gnd 7.36fF $ **FLOATING
C266 a_17685_3840.n35 gnd 7.36fF $ **FLOATING
C267 a_17685_3840.n36 gnd 7.36fF $ **FLOATING
C268 a_17685_3840.n37 gnd 7.36fF $ **FLOATING
C269 a_17685_3840.n38 gnd 7.36fF $ **FLOATING
C270 a_17685_3840.n39 gnd 7.36fF $ **FLOATING
C271 a_17685_3840.n40 gnd 7.36fF $ **FLOATING
C272 a_17685_3840.n41 gnd 7.36fF $ **FLOATING
C273 a_17685_3840.t52 gnd 2.78fF $ **FLOATING
C274 a_17685_3840.n42 gnd 6.20fF $ **FLOATING
C275 a_17685_3840.t39 gnd 3.73fF $ **FLOATING
C276 a_17685_3840.n43 gnd 7.69fF $ **FLOATING
C277 a_17685_3840.t45 gnd 2.78fF $ **FLOATING
C278 a_17685_3840.t37 gnd 2.78fF $ **FLOATING
C279 a_17685_3840.t30 gnd 2.78fF $ **FLOATING
C280 a_17685_3840.t32 gnd 2.78fF $ **FLOATING
C281 a_17685_3840.t23 gnd 2.78fF $ **FLOATING
C282 a_17685_3840.t17 gnd 2.78fF $ **FLOATING
C283 a_17685_3840.t40 gnd 2.78fF $ **FLOATING
C284 a_17685_3840.t34 gnd 2.78fF $ **FLOATING
C285 a_17685_3840.t25 gnd 2.78fF $ **FLOATING
C286 a_17685_3840.t19 gnd 2.78fF $ **FLOATING
C287 a_17685_3840.t59 gnd 6.42fF $ **FLOATING
C288 a_17685_3840.n44 gnd 11.34fF $ **FLOATING
C289 a_17685_3840.n45 gnd 7.38fF $ **FLOATING
C290 a_17685_3840.n46 gnd 7.38fF $ **FLOATING
C291 a_17685_3840.n47 gnd 7.38fF $ **FLOATING
C292 a_17685_3840.n48 gnd 7.38fF $ **FLOATING
C293 a_17685_3840.n49 gnd 7.38fF $ **FLOATING
C294 a_17685_3840.n50 gnd 7.38fF $ **FLOATING
C295 a_17685_3840.n51 gnd 7.38fF $ **FLOATING
C296 a_17685_3840.n52 gnd 7.38fF $ **FLOATING
C297 a_17685_3840.n53 gnd 6.24fF $ **FLOATING
C298 a_17685_3840.t26 gnd 3.73fF $ **FLOATING
C299 a_17685_3840.n54 gnd 5.42fF $ **FLOATING
C300 a_17685_3840.n55 gnd 6.23fF $ **FLOATING
C301 a_17685_3840.n56 gnd 3.39fF $ **FLOATING
C302 a_17685_3840.n61 gnd 2.24fF $ **FLOATING
C303 a_25099_11445.n0 gnd 4.85fF $ **FLOATING
C304 a_25099_11445.t40 gnd 9.08fF $ **FLOATING
C305 a_25099_11445.t15 gnd 10.03fF $ **FLOATING
C306 a_25099_11445.n3 gnd 2.56fF $ **FLOATING
C307 a_25099_11445.t53 gnd 8.63fF $ **FLOATING
C308 a_25099_11445.n4 gnd 7.06fF $ **FLOATING
C309 CLK_BY_4_IPH.t0 gnd 8.55fF
C310 CLK_BY_4_IPH.n3 gnd 30.42fF $ **FLOATING
C311 a_26036_4988.n0 gnd 9.29fF $ **FLOATING
C312 a_26036_4988.n1 gnd 4.19fF $ **FLOATING
C313 a_26036_4988.t20 gnd 9.20fF $ **FLOATING
C314 a_26036_4988.t44 gnd 6.43fF $ **FLOATING
C315 a_26036_4988.t16 gnd 5.98fF $ **FLOATING
C316 vbiasr.t20 gnd 33.23fF
C317 vbiasr.n16 gnd 125.06fF $ **FLOATING
C318 vbiasr.n27 gnd 4.08fF $ **FLOATING
C319 vbiasr.n28 gnd 4.05fF $ **FLOATING
C320 vbiasr.n39 gnd 3.07fF $ **FLOATING
C321 Fvco_By4_QPH.n1 gnd 11.39fF $ **FLOATING
C322 Fvco_By4_QPH.n3 gnd 2.48fF $ **FLOATING
C323 Fvco_By4_QPH.n4 gnd 2.45fF $ **FLOATING
C324 Fvco_By4_QPH.n5 gnd 5.17fF $ **FLOATING
C325 Fvco_By4_QPH.n7 gnd 5.63fF $ **FLOATING
C326 a_49874_4150.n0 gnd 4.09fF $ **FLOATING
C327 a_49874_4150.t6 gnd 2.43fF $ **FLOATING
C328 a_49874_4150.t12 gnd 2.48fF $ **FLOATING
C329 a_49874_4150.t9 gnd 2.26fF $ **FLOATING
C330 a_14188_14050.n0 gnd 9.38fF $ **FLOATING
C331 a_14188_14050.t39 gnd 4.60fF $ **FLOATING
C332 a_14188_14050.t31 gnd 20.11fF $ **FLOATING
C333 a_14188_14050.n3 gnd 3.53fF $ **FLOATING
C334 a_14188_14050.t12 gnd 10.19fF $ **FLOATING
C335 a_14188_14050.n4 gnd 10.20fF $ **FLOATING
C336 a_26690_784.n0 gnd 3.33fF $ **FLOATING
C337 a_23414_5032.n0 gnd 7.44fF $ **FLOATING
C338 a_23414_5032.t14 gnd 13.39fF $ **FLOATING
C339 a_23414_5032.n4 gnd 2.40fF $ **FLOATING
C340 a_23414_5032.t2 gnd 6.75fF $ **FLOATING
C341 a_23414_5032.n5 gnd 5.65fF $ **FLOATING
C342 a_26368_16652.n0 gnd 4.19fF $ **FLOATING
C343 a_26368_16652.t52 gnd 11.90fF $ **FLOATING
C344 a_26368_16652.t39 gnd 9.00fF $ **FLOATING
C345 a_26368_16652.t24 gnd 6.01fF $ **FLOATING
C346 a_26368_16652.n3 gnd 4.12fF $ **FLOATING
C347 Fvco_By4_QPH_bar.n0 gnd 21.37fF $ **FLOATING
C348 Fvco_By4_QPH_bar.n2 gnd 3.86fF $ **FLOATING
C349 Fvco_By4_QPH_bar.n3 gnd 3.48fF $ **FLOATING
C350 Fvco_By4_QPH_bar.n5 gnd 7.86fF $ **FLOATING
