* NGSPICE file created from a.ext - technology: sky130A

X0 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X2 a_28994_17218# a_26368_16652.t2 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X3 a_26690_784.t0 a_23414_5032.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X4 vdd vdd vbiasr.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X5 vinit.t39 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X6 vdd Vso1b a_4226_11420# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X7 vdd reset a_64884_26512# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X8 a_28220_17218# a_26368_16652.t3 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X9 a_29510_17218# a_26368_16652.t4 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X10 a_23403_5596# a_14188_14050.t2 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X11 a_22629_5596# a_14188_14050.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X12 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X13 a_50320_14126# Fvco_By4_QPH.t4 a_55602_11692# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=1.98421e+11p ps=1.49053e+06u w=1e+06u l=150000u
X14 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X15 a_65470_24957# a_64225_24908.t2 a_65009_25170# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.792e+11p pd=1.62e+06u as=2.41013e+11p ps=1.515e+06u w=840000u l=150000u
X16 a_64506_25292# a_33900_31430.t5 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=9.09625e+10p ps=656213u w=420000u l=150000u
X17 a_29510_17218# a_26368_16652.t5 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X18 a_28994_5597# a_26036_4988.t2 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X19 a_22887_5596# a_14188_14050.t4 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X20 a_9354_33563# a_33804_31120.t5 vctrl gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=3.012e+11p ps=2.62e+06u w=1e+06u l=150000u
X21 a_63262_26170# a_61865_26121.t2 a_63110_26170# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.45098e+11p ps=990566u w=420000u l=150000u
X22 a_26847_11500# a_25099_11445.t2 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X23 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X24 a_24177_5596# a_14188_14050.t5 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X25 gnd a_17685_3840.t13 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X26 a_22629_11500# a_14266_8900.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X27 gnd a_17685_3840.t14 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X28 vbiasob.t1 vbiasob.t0 a_54432_7362.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X29 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X30 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X31 a_28736_5597# a_26036_4988.t3 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X32 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X33 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X34 a_26847_11500# a_25099_11445.t3 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X35 a_29510_5597# a_26036_4988.t4 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X36 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X37 gnd Vso3b a_8744_13422# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X38 gnd a_17685_3840.t15 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X39 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X40 a_65009_25170# a_64835_25020# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.41013e+11p pd=1.515e+06u as=1.81925e+11p ps=1.31243e+06u w=840000u l=150000u
X41 gnd Vso5b a_8748_12270# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X42 a_26847_11500# a_25099_11445.t4 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X43 a_23919_5596# a_14188_14050.t6 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X44 a_28994_5597# a_26036_4988.t5 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X45 vdd vdd vbiasr.t18 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X46 a_52052_20860.t18 a_56334_20860.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X47 a_26847_11500# a_25099_11445.t5 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X48 a_23156_5032.t6 a_14188_14050.t7 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X49 a_28736_17218# a_26368_16652.t6 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X50 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X51 a_64394_24908# a_64225_24908.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X52 a_25299_17217# a_23436_16644.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X53 gnd gnd vbiasr.t39 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X54 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X55 a_26847_17217# a_23436_16644.t3 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X56 a_28736_17218# a_26368_16652.t7 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X57 a_25815_5596# a_23414_5032.t3 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X58 a_51276_14152# Fvco_By4_QPH.t5 a_51636_13108# gnd sky130_fd_pr__nfet_01v8 ad=2.07143e+11p pd=1.67714e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X59 gnd a_17685_3840.t16 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X60 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X61 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X62 a_23145_5596# a_14188_14050.t8 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X63 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X64 vdd a_63110_26170# a_62307_26207# vdd sky130_fd_pr__pfet_01v8_hvt ad=2.72887e+11p pd=1.96864e+06u as=1.764e+11p ps=1.54e+06u w=1.26e+06u l=150000u
X65 a_26331_11500# a_25099_11445.t6 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X66 a_28478_5597# a_26036_4988.t6 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X67 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X68 vdd reset a_62146_26505# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X69 a_29252_5597# a_26036_4988.t7 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X70 vdd Fvco a_4288_11534# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X71 a_25778_4988.t6 a_23414_5032.t4 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X72 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X73 a_26331_11500# a_25099_11445.t7 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X74 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X75 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X76 gnd a_63282_26362# a_63262_26170# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=4.41e+10p ps=630000u w=420000u l=150000u
X77 gnd a_17685_3840.t17 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X78 a_23145_17217# a_22429_17162.t2 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X79 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X80 a_28220_17218# a_26368_16652.t8 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X81 a_23145_17217# a_22429_17162.t3 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X82 a_52052_20860.t8 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X83 a_56602_11692# vbiasob.t3 a_56272_15934.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=2e+06u
X84 a_27962_5597# a_26036_4988.t8 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X85 a_26331_17217# a_23436_16644.t4 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X86 a_28220_17218# a_26368_16652.t9 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X87 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X88 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X89 a_63420_26170# reset gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=9.24629e+10p ps=686014u w=420000u l=150000u
X90 a_25557_11500# a_25099_11445.t8 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X91 a_25557_5596# a_23414_5032.t5 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X92 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X93 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X94 a_49916_3664.t0 a_49858_3690.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.81792e+11p ps=2.09071e+06u w=1.28e+06u l=8e+06u
X95 a_22887_5596# a_14188_14050.t9 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X96 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X97 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X98 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X99 a_49858_3690.t1 a_49858_3690.t0 a_54934_4354# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.856e+11p ps=1.57e+06u w=1.28e+06u l=8e+06u
X100 a_23661_5596# a_14188_14050.t10 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X101 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X102 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X103 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X104 a_26847_5596# a_23414_5032.t6 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X105 a_28578_5014.t6 a_26036_4988.t9 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X106 a_51516_3690.t2 a_51516_3690.t1 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.59518e+11p ps=2.5936e+06u w=1.66e+06u l=4e+06u
X107 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X108 a_62265_26233# reset gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=9.24629e+10p ps=686014u w=420000u l=150000u
X109 a_28220_5597# a_26036_4988.t10 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X110 gnd a_17685_3840.t18 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X111 a_24177_11500# a_14266_8900.t3 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X112 a_50583_13108.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X113 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X114 a_25557_11500# a_25099_11445.t9 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X115 a_52052_20860.t17 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X116 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X117 a_23403_5596# a_14188_14050.t11 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X118 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X119 vdd a_66604_26416# Fvco_By4_QPH_bar.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=2.72887e+11p pd=1.96864e+06u as=0p ps=0u w=1.26e+06u l=150000u
X120 a_29252_11501# a_27762_11446.t2 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X121 a_25557_11500# a_25099_11445.t10 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X122 a_25299_5596# a_23414_5032.t7 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X123 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X124 a_28994_5597# a_26036_4988.t11 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X125 vdd vdd vinit.t19 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X126 a_25557_11500# a_25099_11445.t11 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X127 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X128 a_65360_26240# a_64772_26128# a_65213_26240# gnd sky130_fd_pr__nfet_01v8 ad=4.935e+10p pd=655000u as=1.2285e+11p ps=1.005e+06u w=420000u l=150000u
X129 vbiasr.t38 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X130 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X131 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X132 a_26589_5596# a_23414_5032.t8 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X133 a_24177_11500# a_14266_8900.t4 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X134 a_44752_16348.t2 a_51138_19904.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X135 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X136 a_25557_17217# a_23436_16644.t5 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X137 a_24177_11500# a_14266_8900.t5 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X138 a_27962_11501# a_27762_11446.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X139 gnd gnd vbiasr.t37 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X140 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X141 a_14832_12082.t0 a_14188_14050.t12 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X142 a_29252_11501# a_27762_11446.t4 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X143 a_56602_11692# a_51636_13108# a_52052_20860.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X144 a_29510_5597# a_26036_4988.t12 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X145 a_24177_11500# a_14266_8900.t6 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X146 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X147 a_33808_31746# a_33900_31430.t6 a_34044_31208# vdd sky130_fd_pr__pfet_01v8 ad=3.78914e+11p pd=2.83143e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X148 a_63282_26362# a_63110_26170# a_63420_26170# gnd sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=4.41e+10p ps=630000u w=420000u l=150000u
X149 a_29252_11501# a_27762_11446.t5 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X150 vdd a_56334_19906# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X151 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X152 a_26073_5596# a_23414_5032.t9 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X153 a_24177_17217# a_22429_17162.t4 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X154 a_29252_11501# a_27762_11446.t6 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X155 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X156 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X157 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X158 a_64884_26512# Fvco_By4_QPH.t6 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=9.09625e+10p ps=656213u w=420000u l=150000u
X159 a_26847_17217# a_23436_16644.t6 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X160 a_23160_10936.t7 a_14266_8900.t7 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X161 gnd Vso7b a_8748_11114# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X162 a_29252_17218# a_26368_16652.t10 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X163 a_23661_11500# a_14266_8900.t8 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X164 a_26847_17217# a_23436_16644.t7 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X165 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X166 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X167 a_62146_26505# a_62307_26207# a_62265_26233# gnd sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=960000u as=4.41e+10p ps=630000u w=420000u l=150000u
X168 a_64066_26111# a_63866_26409# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.54e+06u as=2.72887e+11p ps=1.96864e+06u w=1.26e+06u l=150000u
X169 a_23661_11500# a_14266_8900.t9 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X170 a_25815_5596# a_23414_5032.t10 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X171 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X172 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X173 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X174 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X175 a_23919_11500# a_14266_8900.t10 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X176 a_26331_5596# a_23414_5032.t11 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X177 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X178 a_55602_11692# a_51041_13108# a_52052_20860.t16 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X179 a_42574_15624# Fvco_By4_QPH_bar.t4 a_42550_16062# vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X180 a_29252_5597# a_26036_4988.t13 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X181 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X182 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X183 vinit.t18 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X184 a_23661_17217# a_22429_17162.t5 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X185 a_26331_17217# a_23436_16644.t8 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X186 a_22887_11500# a_14266_8900.t11 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X187 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X188 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X189 a_28438_10874.t6 a_27762_11446.t7 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X190 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X191 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X192 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X193 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X194 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X195 gnd gnd vinit.t38 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X196 gnd a_17685_3840.t19 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X197 a_26331_17217# a_23436_16644.t9 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X198 a_23919_11500# a_14266_8900.t12 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X199 gnd a_17685_3840.t20 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X200 a_28438_10874.t5 a_27762_11446.t8 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X201 a_25557_5596# a_23414_5032.t12 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X202 vinit.t17 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X203 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X204 gnd a_63110_26170# a_62307_26207# gnd sky130_fd_pr__nfet_01v8 ad=1.84926e+11p pd=1.37203e+06u as=1.176e+11p ps=1.12e+06u w=840000u l=150000u
X205 a_23919_11500# a_14266_8900.t13 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X206 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X207 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X208 a_23919_11500# a_14266_8900.t14 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X209 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X210 gnd a_17685_3840.t21 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X211 a_22887_11500# a_14266_8900.t15 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X212 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X213 a_14910_6932.t0 a_14266_8900.t16 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X214 vbiasr.t36 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X215 a_28622_16652# a_26368_16652.t11 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X216 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X217 gnd Vso4b a_8740_12844# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X218 a_4314_11564# a_4288_11534# a_4314_11468# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X219 a_23919_17217# a_22429_17162.t6 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X220 a_22887_11500# a_14266_8900.t17 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X221 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X222 gnd a_17685_3840.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X223 gnd a_17685_3840.t23 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X224 vdd a_4288_11918# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X225 a_23403_11500# a_14266_8900.t18 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X226 a_22887_11500# a_14266_8900.t19 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X227 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X228 a_64835_25020# a_64225_24908.t4 a_64506_25292# gnd sky130_fd_pr__nfet_01v8 ad=1.2285e+11p pd=1.005e+06u as=1.134e+11p ps=960000u w=420000u l=150000u
X229 a_64066_26111# a_63866_26409# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.12e+06u as=1.84926e+11p ps=1.37203e+06u w=840000u l=150000u
X230 a_65213_26240# a_64603_26128.t2 a_64884_26512# gnd sky130_fd_pr__nfet_01v8 ad=1.2285e+11p pd=1.005e+06u as=1.134e+11p ps=960000u w=420000u l=150000u
X231 a_23403_11500# a_14266_8900.t20 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X232 a_26016_10878.t6 a_25099_11445.t12 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X233 a_25299_5596# a_23414_5032.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X234 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X235 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X236 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X237 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X238 a_22887_17217# a_22429_17162.t7 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X239 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X240 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X241 a_28622_16652# a_26368_16652.t12 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X242 a_25557_17217# a_23436_16644.t10 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X243 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X244 gnd a_17685_3840.t24 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X245 a_25557_17217# a_23436_16644.t11 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X246 a_26073_11500# a_25099_11445.t13 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X247 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X248 a_23403_17217# a_22429_17162.t8 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X249 a_64835_25020# reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=7.63e+10p pd=923333u as=9.09625e+10p ps=656213u w=420000u l=150000u
X250 a_22629_11500# a_14266_8900.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X251 a_62631_26505# a_61865_26121.t3 a_62475_26233# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.41e+10p pd=630000u as=7.63e+10p ps=923333u w=420000u l=150000u
X252 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X253 a_77280_24640.t1 a_77254_23336.t4 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X254 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X255 a_65059_25020# a_65009_25170# a_64982_25020# gnd sky130_fd_pr__nfet_01v8 ad=5.775e+10p pd=695000u as=4.935e+10p ps=655000u w=420000u l=150000u
X256 a_24177_17217# a_22429_17162.t9 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X257 vbiasr.t17 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X258 vbiasr.t35 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X259 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X260 a_24177_17217# a_22429_17162.t10 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X261 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X262 a_29252_17218# a_26368_16652.t13 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X263 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X264 Vso1b a_24410_25128.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X265 a_28478_11501# a_27762_11446.t9 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X266 a_49916_3664.t2 a_49916_3664.t1 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16577e+11p ps=1.56241e+06u w=1e+06u l=2e+07u
X267 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X268 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X269 vinit.t37 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X270 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X271 a_29252_17218# a_26368_16652.t14 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X272 a_22629_11500# a_14266_8900.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X273 a_23308_802.t1 a_22429_17162.t11 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X274 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X275 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X276 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X277 a_26368_16652.t1 a_23436_16644.t12 a_26110_16652# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X278 a_28478_11501# a_27762_11446.t10 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X279 a_24177_5596# a_14188_14050.t13 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X280 a_57710_5326.t0 a_51516_3690.t4 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.72513e+11p ps=2.68735e+06u w=1.72e+06u l=4e+06u
X281 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.2015e+11p pd=1.63337e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X282 a_22629_11500# a_14266_8900.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X283 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X284 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X285 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X286 vdd Fvco a_61865_26121.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38609e+11p pd=999944u as=0p ps=0u w=640000u l=150000u
X287 gnd a_64066_26111# a_64603_26128.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=0p ps=0u w=420000u l=150000u
X288 a_22629_11500# a_14266_8900.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X289 a_23661_17217# a_22429_17162.t12 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X290 gnd Vso1b a_8744_9386# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X291 a_28478_17218# a_26368_16652.t15 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X292 a_57710_5326.t4 a_57710_5326.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.60449e+11p ps=4.9001e+06u w=3e+06u l=1e+06u
X293 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X294 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X295 vdd a_65470_24957# a_66226_25196# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38609e+11p pd=999944u as=1.696e+11p ps=1.81e+06u w=640000u l=150000u
X296 a_22629_17217# a_22429_17162.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X297 a_23661_17217# a_22429_17162.t14 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X298 a_26036_4988.t0 a_23414_5032.t14 a_17685_3840.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X299 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X300 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X301 vdd a_4226_11420# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X302 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X303 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X304 vbiasr.t16 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X305 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X306 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X307 vdd a_4226_12188# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X308 a_25815_11500# a_25099_11445.t14 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X309 a_32948_24994.t0 a_27762_11446.t11 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X310 Vso2b a_28790_25040.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X311 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X312 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X313 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X314 vdd vdd vinit.t16 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X315 a_33804_31120.t3 a_66226_25196# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.84926e+11p ps=1.37203e+06u w=840000u l=150000u
X316 a_28478_17218# a_26368_16652.t16 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X317 vdd a_66020_26369# a_65978_26545# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=4.41e+10p ps=630000u w=420000u l=150000u
X318 a_28622_16652# a_26368_16652.t17 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X319 a_23145_5596# a_14188_14050.t14 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X320 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X321 a_23919_17217# a_22429_17162.t15 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X322 a_65780_24957# reset gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=9.24629e+10p ps=686014u w=420000u l=150000u
X323 gnd a_17685_3840.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X324 a_28622_16652# a_26368_16652.t18 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X325 a_62034_26121# a_61865_26121.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X326 a_23919_17217# a_22429_17162.t16 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X327 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X328 a_14910_6932.t1 a_14266_8900.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X329 gnd a_17685_3840.t26 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X330 a_52052_20860.t6 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X331 gnd a_17685_3840.t27 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X332 vdd vdd vinit.t15 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X333 a_51276_14152# a_51334_14126# a_33808_31746# gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=3.78571e+11p ps=2.99714e+06u w=2e+06u l=1e+06u
X334 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X335 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X336 vdd Vso6b a_4226_11804# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X337 a_22887_17217# a_22429_17162.t17 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X338 a_29510_11501# a_27762_11446.t12 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X339 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X340 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X341 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X342 a_64835_25020# a_64394_24908# a_64506_25292# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.63e+10p pd=923333u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X343 a_27962_5597# a_26036_4988.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X344 a_22887_17217# a_22429_17162.t18 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X345 vbiasr.t15 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X346 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X347 a_56602_11692# a_51636_13108# a_52052_20860.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X348 vdd a_50032_16080.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X349 a_23403_17217# a_22429_17162.t19 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X350 a_23661_5596# a_14188_14050.t15 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X351 a_22887_5596# a_14188_14050.t16 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X352 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X353 a_50511_16072.t5 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X354 a_64625_25020# reset gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=9.24629e+10p ps=686014u w=420000u l=150000u
X355 a_23403_17217# a_22429_17162.t20 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X356 a_23919_5596# a_14188_14050.t17 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X357 vdd a_51138_19904.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X358 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X359 a_62622_26233# a_62034_26121# a_62475_26233# gnd sky130_fd_pr__nfet_01v8 ad=4.935e+10p pd=655000u as=1.2285e+11p ps=1.005e+06u w=420000u l=150000u
X360 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X361 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X362 vdd a_62307_26207# a_64225_24908.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38609e+11p pd=999944u as=0p ps=0u w=640000u l=150000u
X363 a_52052_20860.t15 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X364 a_50583_13108.t0 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X365 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X366 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X367 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X368 a_27962_11501# a_27762_11446.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X369 Vso4b a_38070_8852.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X370 a_52052_20224# a_56272_15934.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X371 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X372 a_14266_8900.t1 a_25099_11445.t15 a_26016_10878.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X373 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X374 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X375 vdd a_65848_26177# Fvco_By4_QPH.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=2.72887e+11p pd=1.96864e+06u as=0p ps=0u w=1.26e+06u l=150000u
X376 a_28994_5597# a_26036_4988.t15 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X377 Vso5b a_14910_6932.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X378 a_26589_11500# a_25099_11445.t16 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X379 a_65642_25149# a_65470_24957# a_65780_24957# gnd sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=4.41e+10p ps=630000u w=420000u l=150000u
X380 a_55602_11692# a_51041_13108# a_52052_20860.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X381 a_26589_11500# a_25099_11445.t17 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X382 a_23919_5596# a_14188_14050.t18 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X383 a_24177_5596# a_14188_14050.t19 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X384 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X385 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X386 a_63282_26362# reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=9.09625e+10p ps=656213u w=420000u l=150000u
X387 gnd a_66020_26369# a_66000_26177# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=4.41e+10p ps=630000u w=420000u l=150000u
X388 a_23160_10936.t6 a_14266_8900.t26 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X389 a_27962_11501# a_27762_11446.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X390 a_56602_11692# a_51636_13108# a_52052_20860.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X391 vinit.t14 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X392 a_27962_11501# a_27762_11446.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X393 a_49858_3690.t2 a_51516_3690.t5 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.59518e+11p ps=2.5936e+06u w=1.66e+06u l=4e+06u
X394 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X395 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X396 a_28478_17218# a_26368_16652.t19 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X397 a_30384_802.t0 a_26036_4988.t16 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X398 a_77598_24640.t1 a_77572_23336.t3 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X399 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X400 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X401 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X402 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X403 a_4314_12044# a_4226_11996# a_4314_11948# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X404 a_26589_17217# a_23436_16644.t13 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X405 a_22629_17217# a_22429_17162.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X406 a_27962_11501# a_27762_11446.t16 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X407 a_28478_17218# a_26368_16652.t20 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X408 a_26073_5596# a_23414_5032.t15 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X409 a_22629_17217# a_22429_17162.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X410 a_23145_11500# a_14266_8900.t27 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X411 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X412 a_23160_10936.t5 a_14266_8900.t28 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X413 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X414 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X415 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X416 a_27962_17218# a_26368_16652.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X417 a_51041_13108# a_50511_16072.t8 a_50583_13108.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X418 a_64506_25292# a_33900_31430.t7 a_64625_25020# gnd sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=960000u as=4.41e+10p ps=630000u w=420000u l=150000u
X419 a_23160_10936.t4 a_14266_8900.t29 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X420 a_28220_11501# a_27762_11446.t17 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X421 a_28578_5014.t5 a_26036_4988.t17 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X422 a_23160_10936.t3 a_14266_8900.t30 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X423 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X424 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X425 a_26847_17217# a_23436_16644.t14 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X426 a_53292_3120# a_49858_3690.t5 vbiasr.t40 gnd sky130_fd_pr__nfet_01v8 ad=7.0035e+11p pd=5.12e+06u as=0p ps=0u w=4.83e+06u l=8e+06u
X427 a_55602_11692# a_51041_13108# a_52052_20860.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X428 a_23403_5596# a_14188_14050.t20 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X429 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X430 vdd vdd vinit.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X431 a_23178_16644# a_22429_17162.t23 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X432 Fvco a_23308_802.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X433 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X434 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X435 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X436 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X437 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X438 a_64772_26128# a_64603_26128.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.696e+11p pd=1.81e+06u as=1.38609e+11p ps=999944u w=640000u l=150000u
X439 gnd a_17685_3840.t28 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X440 gnd a_17685_3840.t29 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X441 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X442 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X443 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X444 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X445 a_28578_5014.t4 a_26036_4988.t18 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X446 gnd Vso2b a_8736_14034# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X447 a_27962_5597# a_26036_4988.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X448 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X449 vinit.t36 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X450 vdd a_4226_11996# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X451 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X452 gnd a_17685_3840.t30 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X453 a_22429_17162.t1 a_26036_4988.t20 a_28578_5014.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X454 a_22629_5596# a_14188_14050.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X455 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X456 a_26016_10878.t5 a_25099_11445.t18 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X457 a_25299_11500# a_25099_11445.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X458 a_29510_5597# a_26036_4988.t21 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X459 a_23403_5596# a_14188_14050.t22 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X460 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X461 a_23661_5596# a_14188_14050.t23 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X462 a_25299_11500# a_25099_11445.t20 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X463 a_23919_5596# a_14188_14050.t24 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X464 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X465 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X466 gnd a_17685_3840.t31 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X467 gnd a_65848_26177# a_66604_26416# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X468 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X469 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X470 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X471 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X472 a_26073_11500# a_25099_11445.t21 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X473 vdd vdd vbiasr.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X474 gnd gnd vbiasr.t34 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X475 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X476 a_25299_17217# a_23436_16644.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X477 Vso7b a_26690_784.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X478 a_30384_802.t1 a_26036_4988.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X479 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X480 a_26016_10878.t4 a_25099_11445.t22 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X481 a_25815_5596# a_23414_5032.t16 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X482 a_28736_5597# a_26036_4988.t23 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X483 a_26016_10878.t3 a_25099_11445.t23 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X484 a_29252_5597# a_26036_4988.t24 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X485 a_29510_5597# a_26036_4988.t25 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X486 a_65213_26240# a_64772_26128# a_64884_26512# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.63e+10p pd=923333u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X487 a_26016_10878.t2 a_25099_11445.t24 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X488 a_66000_26177# a_64603_26128.t4 a_65848_26177# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.45098e+11p ps=990566u w=420000u l=150000u
X489 gnd a_17685_3840.t32 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X490 a_26073_11500# a_25099_11445.t25 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X491 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X492 a_56602_11692# Fvco_By4_QPH_bar.t5 a_50320_14126# gnd sky130_fd_pr__nfet_01v8 ad=1.98421e+11p pd=1.49053e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X493 a_23156_5032.t5 a_14188_14050.t25 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X494 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X495 gnd a_17685_3840.t33 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X496 a_46856_21176.t1 a_51138_21494.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X497 gnd a_17685_3840.t34 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X498 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X499 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X500 a_26110_16652# a_23436_16644.t16 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X501 a_25557_17217# a_23436_16644.t17 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X502 a_26073_11500# a_25099_11445.t26 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X503 a_26589_17217# a_23436_16644.t18 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X504 a_77280_24640.t2 a_77254_23336.t3 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X505 a_26073_11500# a_25099_11445.t27 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X506 gnd gnd vinit.t35 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X507 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X508 a_26589_17217# a_23436_16644.t19 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X509 a_25815_5596# a_23414_5032.t17 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X510 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X511 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X512 gnd a_65848_26177# Fvco_By4_QPH.t3 gnd sky130_fd_pr__nfet_01v8 ad=1.84926e+11p pd=1.37203e+06u as=0p ps=0u w=840000u l=150000u
X513 a_27962_17218# a_26368_16652.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X514 a_25557_5596# a_23414_5032.t18 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X515 a_42574_15624# vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=4e+06u
X516 gnd a_56334_20860.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X517 a_26073_5596# a_23414_5032.t19 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X518 a_28478_5597# a_26036_4988.t26 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X519 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X520 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X521 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X522 gnd gnd vbiasr.t33 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X523 a_29252_5597# a_26036_4988.t27 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X524 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X525 a_26073_17217# a_23436_16644.t20 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X526 a_24177_17217# a_22429_17162.t24 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X527 a_27962_17218# a_26368_16652.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X528 a_25778_4988.t5 a_23414_5032.t20 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X529 gnd a_17685_3840.t35 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X530 a_26331_11500# a_25099_11445.t28 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X531 gnd gnd vinit.t34 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X532 a_28578_5014.t3 a_26036_4988.t28 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X533 vdd Vso3b a_4288_12110# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X534 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X535 vdd Vso5b a_4288_11918# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X536 a_23178_16644# a_22429_17162.t25 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X537 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X538 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X539 a_34044_31208# a_33804_31120.t6 a_33808_31746# gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=1.89286e+11p ps=1.49857e+06u w=1e+06u l=150000u
X540 Vso3b a_32948_24994.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X541 a_25815_11500# a_25099_11445.t29 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X542 a_23403_5596# a_14188_14050.t26 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X543 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X544 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X545 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X546 a_23178_16644# a_22429_17162.t26 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X547 a_25557_5596# a_23414_5032.t21 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X548 a_23504_23306# vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X549 a_25299_5596# a_23414_5032.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X550 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X551 a_33808_31746# a_33900_31430.t8 a_9354_33563# gnd sky130_fd_pr__nfet_01v8 ad=1.89286e+11p pd=1.49857e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X552 vdd a_65848_26177# a_66020_26369# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=5.88e+10p ps=700000u w=420000u l=150000u
X553 a_51636_13108# a_50511_16072.t9 a_46856_19268.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X554 a_77280_24640.t0 a_33900_31430.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X555 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X556 vdd a_63282_26362# a_63240_26538# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=4.41e+10p ps=630000u w=420000u l=150000u
X557 a_26847_5596# a_23414_5032.t23 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X558 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X559 a_25815_11500# a_25099_11445.t30 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X560 gnd gnd vbiasr.t32 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X561 a_45810_16322# Fvco_By4_QPH.t7 a_47968_16078# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X562 a_28220_5597# a_26036_4988.t29 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X563 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X564 vdd Vso7b a_4226_11612# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X565 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X566 a_29510_11501# a_27762_11446.t18 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X567 a_25815_11500# a_25099_11445.t31 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X568 a_29510_5597# a_26036_4988.t30 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X569 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X570 vinit.t12 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X571 a_25815_11500# a_25099_11445.t32 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X572 a_47968_16078# Fvco_By4_QPH_bar.t6 a_44810_16322# vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X573 a_65213_26240# reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=7.63e+10p pd=923333u as=9.09625e+10p ps=656213u w=420000u l=150000u
X574 a_25299_5596# a_23414_5032.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X575 vdd vdd vbiasr.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X576 vbiasot.t0 a_51516_3690.t6 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16952e+11p ps=843703u w=540000u l=8e+06u
X577 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X578 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X579 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X580 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X581 Vso3b a_32948_24994.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X582 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X583 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X584 vdd Vso7b a_4288_11726# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X585 a_25815_17217# a_23436_16644.t21 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X586 a_25299_17217# a_23436_16644.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X587 a_26589_5596# a_23414_5032.t25 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X588 a_23919_17217# a_22429_17162.t27 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X589 a_9354_33563# a_33804_31120.t7 a_33808_31746# vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.78914e+11p ps=2.83143e+06u w=2e+06u l=150000u
X590 a_25299_17217# a_23436_16644.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X591 a_29510_11501# a_27762_11446.t19 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X592 a_25815_5596# a_23414_5032.t26 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X593 a_29510_11501# a_27762_11446.t20 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X594 Fvco a_23308_802.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X595 a_25099_11445.t0 a_27762_11446.t21 a_28438_10874.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X596 a_28790_25040.t0 a_26368_16652.t24 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X597 a_22887_17217# a_22429_17162.t28 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X598 a_29510_11501# a_27762_11446.t22 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X599 a_29252_5597# a_26036_4988.t31 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X600 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X601 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X602 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X603 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X604 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X605 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X606 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X607 a_26110_16652# a_23436_16644.t24 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X608 vdd vdd vbiasr.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X609 Vso5b a_14910_6932.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X610 a_23436_16644.t1 a_22429_17162.t29 a_17685_3840.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X611 vinit.t11 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X612 a_29510_17218# a_26368_16652.t25 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X613 Vso7b a_26690_784.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X614 a_26110_16652# a_23436_16644.t25 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X615 a_77598_24640.t2 a_77572_23336.t2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X616 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X617 vdd a_65848_26177# a_66604_26416# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38609e+11p pd=999944u as=1.696e+11p ps=1.81e+06u w=640000u l=150000u
X618 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X619 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X620 a_23661_11500# a_14266_8900.t31 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X621 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X622 a_26073_17217# a_23436_16644.t26 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X623 a_25557_5596# a_23414_5032.t27 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X624 vdd Vso8b a_4288_11534# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X625 a_26331_5596# a_23414_5032.t28 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X626 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X627 gnd a_17685_3840.t36 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X628 a_26073_17217# a_23436_16644.t27 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X629 gnd a_17685_3840.t37 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X630 a_50262_14152# Fvco_By4_QPH.t8 a_51041_13108# gnd sky130_fd_pr__nfet_01v8 ad=2.07143e+11p pd=1.67714e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X631 a_47968_16078# a_42550_16062# a_50511_16072.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X632 a_23145_11500# a_14266_8900.t32 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X633 vdd Fvco a_4226_11420# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X634 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X635 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X636 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X637 a_45810_16322# vbiasbuffer.t3 a_51826_16054.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=1e+06u
X638 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X639 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X640 vinit.t33 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X641 a_28220_11501# a_27762_11446.t23 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X642 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X643 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X644 gnd reset a_62699_26233# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=5.775e+10p ps=695000u w=420000u l=150000u
X645 vbiasr.t11 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X646 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.0821e+12p pd=2.28671e+07u as=3.0821e+12p ps=2.28671e+07u w=1.4e+07u l=1e+06u
X647 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X648 vdd vdd vinit.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X649 vdd vdd vbiasr.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X650 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X651 a_28438_10874.t4 a_27762_11446.t24 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X652 a_43010_16058# Fvco_By4_QPH.t9 a_42574_15624# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X653 a_25299_5596# a_23414_5032.t29 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X654 a_28994_11501# a_27762_11446.t25 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X655 vinit.t32 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X656 a_23145_11500# a_14266_8900.t33 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X657 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X658 a_22629_17217# a_22429_17162.t30 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X659 a_28994_11501# a_27762_11446.t26 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X660 a_50112_7696# a_54432_7362.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X661 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X662 a_23145_11500# a_14266_8900.t34 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X663 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X664 a_28220_11501# a_27762_11446.t27 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X665 a_23145_11500# a_14266_8900.t35 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X666 a_50511_16072.t4 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X667 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X668 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X669 a_28220_11501# a_27762_11446.t28 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X670 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X671 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X672 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X673 a_23145_17217# a_22429_17162.t31 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X674 a_28994_17218# a_26368_16652.t26 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X675 a_28220_11501# a_27762_11446.t29 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X676 a_42782_16060# vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=4e+06u
X677 a_53292_2532# a_49858_3690.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=2.175e+11p pd=1.79e+06u as=3.30225e+11p ps=2.45005e+06u w=1.5e+06u l=8e+06u
X678 vdd a_51138_19904.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X679 a_77598_24640.t0 a_33804_31120.t4 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X680 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X681 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X682 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X683 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X684 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X685 a_25815_17217# a_23436_16644.t28 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X686 a_23403_11500# a_14266_8900.t36 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X687 a_65848_26177# a_64603_26128.t5 a_65387_26390# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.792e+11p pd=1.62e+06u as=2.41013e+11p ps=1.515e+06u w=840000u l=150000u
X688 a_28220_17218# a_26368_16652.t27 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X689 vdd a_63866_26409# a_64066_26111# vdd sky130_fd_pr__pfet_01v8_hvt ad=2.72887e+11p pd=1.96864e+06u as=1.764e+11p ps=1.54e+06u w=1.26e+06u l=150000u
X690 a_25815_17217# a_23436_16644.t29 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X691 vbiasr.t31 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X692 vctrl a_33900_31430.t9 a_34044_31208# gnd sky130_fd_pr__nfet_01v8 ad=3.012e+11p pd=2.62e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X693 a_52052_20224# a_56334_19906# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X694 a_28994_17218# a_26368_16652.t28 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X695 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X696 a_24177_5596# a_14188_14050.t27 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X697 a_42550_16062# Fvco_By4_QPH.t10 a_42574_15624# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X698 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X699 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X700 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X701 Fvco_By4_QPH_bar.t3 a_66604_26416# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.84926e+11p ps=1.37203e+06u w=840000u l=150000u
X702 a_23436_16644.t0 a_22429_17162.t32 a_23178_16644# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X703 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X704 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X705 a_29510_17218# a_26368_16652.t29 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X706 a_22629_5596# a_14188_14050.t28 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X707 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X708 Vso6b a_14832_12082.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X709 a_28736_11501# a_27762_11446.t30 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X710 gnd a_17685_3840.t38 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X711 gnd gnd vinit.t31 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X712 a_4314_11660# a_4226_11612# a_4314_11564# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X713 a_29510_17218# a_26368_16652.t30 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X714 gnd a_17685_3840.t39 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X715 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X716 a_65387_26390# a_65213_26240# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.41013e+11p pd=1.515e+06u as=1.81925e+11p ps=1.31243e+06u w=840000u l=150000u
X717 a_28736_11501# a_27762_11446.t31 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X718 a_23919_5596# a_14188_14050.t29 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X719 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X720 vinit.t9 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X721 a_28478_11501# a_27762_11446.t32 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X722 a_65848_26177# a_64772_26128# a_65387_26390# gnd sky130_fd_pr__nfet_01v8 ad=2.21102e+11p pd=1.50943e+06u as=1.264e+11p ps=1.035e+06u w=640000u l=150000u
X723 a_24177_5596# a_14188_14050.t30 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X724 a_23414_5032.t1 a_14188_14050.t31 a_17685_3840.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X725 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X726 a_28736_17218# a_26368_16652.t31 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X727 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X728 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X729 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X730 gnd a_17685_3840.t40 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X731 a_28736_5597# a_26036_4988.t32 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X732 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X733 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X734 gnd a_17685_3840.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X735 gnd a_17685_3840.t42 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X736 gnd a_63866_26409# a_64066_26111# gnd sky130_fd_pr__nfet_01v8 ad=1.84926e+11p pd=1.37203e+06u as=1.176e+11p ps=1.12e+06u w=840000u l=150000u
X737 vdd a_65009_25170# a_64991_25292# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=4.41e+10p ps=630000u w=420000u l=150000u
X738 a_26331_11500# a_25099_11445.t33 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X739 a_23156_5032.t4 a_14188_14050.t32 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X740 a_77572_23336.t5 a_77254_23336.t0 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X741 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X742 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X743 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X744 vinit.t30 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X745 a_28736_17218# a_26368_16652.t32 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X746 a_27962_5597# a_26036_4988.t33 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X747 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X748 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X749 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X750 a_4314_11756# a_4288_11726# a_4314_11660# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X751 a_28478_5597# a_26036_4988.t34 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X752 a_23145_5596# a_14188_14050.t33 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X753 a_33804_31120.t1 a_66226_25196# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.72887e+11p ps=1.96864e+06u w=1.26e+06u l=150000u
X754 a_26331_11500# a_25099_11445.t34 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X755 a_23661_5596# a_14188_14050.t34 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X756 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X757 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X758 a_25778_4988.t4 a_23414_5032.t30 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X759 vbiasr.t9 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X760 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X761 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X762 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X763 a_65387_26390# a_65213_26240# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.264e+11p pd=1.035e+06u as=1.40896e+11p ps=1.04535e+06u w=640000u l=150000u
X764 a_28994_17218# a_26368_16652.t33 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X765 a_26331_11500# a_25099_11445.t35 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X766 a_28578_5014.t2 a_26036_4988.t35 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X767 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X768 a_23145_17217# a_22429_17162.t33 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X769 a_23308_802.t0 a_22429_17162.t34 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X770 a_28994_17218# a_26368_16652.t34 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X771 a_26331_11500# a_25099_11445.t36 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X772 a_23145_17217# a_22429_17162.t35 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X773 a_51516_3690.t3 a_49916_3664.t3 a_49858_3690.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.28e+06u l=8e+06u
X774 a_42782_16060# Fvco_By4_QPH_bar.t7 a_43010_16058# vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X775 a_27962_5597# a_26036_4988.t36 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X776 a_28220_17218# a_26368_16652.t35 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X777 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X778 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X779 a_26331_17217# a_23436_16644.t30 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X780 a_23403_5596# a_14188_14050.t35 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X781 a_23178_16644# a_22429_17162.t36 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X782 a_28220_17218# a_26368_16652.t36 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X783 a_51516_3690.t0 a_49858_3690.t7 a_54950_3120# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.0035e+11p ps=5.12e+06u w=4.83e+06u l=8e+06u
X784 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X785 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X786 a_62307_26207# a_63110_26170# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.12e+06u as=1.84926e+11p ps=1.37203e+06u w=840000u l=150000u
X787 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X788 a_22887_5596# a_14188_14050.t36 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X789 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X790 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X791 a_62475_26233# reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=7.63e+10p pd=923333u as=9.09625e+10p ps=656213u w=420000u l=150000u
X792 a_65978_26545# a_64772_26128# a_65848_26177# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.41e+10p pd=630000u as=8.96e+10p ps=810000u w=420000u l=150000u
X793 gnd a_17685_3840.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X794 a_23661_5596# a_14188_14050.t37 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X795 a_54950_3120# a_49858_3690.t8 a_53292_3120# gnd sky130_fd_pr__nfet_01v8 ad=7.0035e+11p pd=5.12e+06u as=7.0035e+11p ps=5.12e+06u w=4.83e+06u l=8e+06u
X796 a_26847_5596# a_23414_5032.t31 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X797 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X798 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X799 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X800 a_64772_26128# a_64603_26128.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X801 vdd Vso8b a_4226_11612# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X802 a_24177_5596# a_14188_14050.t38 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X803 a_28220_5597# a_26036_4988.t37 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X804 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X805 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X806 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X807 vbiasr.t8 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X808 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X809 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X810 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X811 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X812 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X813 vbiasr.t30 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X814 a_46856_19268.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X815 a_23414_5032.t0 a_14188_14050.t39 a_23156_5032.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X816 a_22629_5596# a_14188_14050.t40 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X817 a_26847_11500# a_25099_11445.t37 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X818 a_29510_5597# a_26036_4988.t38 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X819 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X820 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X821 vdd Vso6b a_4288_11726# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X822 a_26073_5596# a_23414_5032.t32 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X823 a_46856_21176.t0 a_51138_20858# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X824 a_26847_11500# a_25099_11445.t38 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X825 a_28994_5597# a_26036_4988.t39 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X826 vbiasot.t2 vbiasot.t1 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=4e+06u
X827 a_26589_11500# a_25099_11445.t39 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X828 a_51826_16054.t1 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X829 gnd a_66226_25196# a_33804_31120.t2 gnd sky130_fd_pr__nfet_01v8 ad=1.84926e+11p pd=1.37203e+06u as=0p ps=0u w=840000u l=150000u
X830 a_26589_5596# a_23414_5032.t33 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X831 a_26036_4988.t1 a_23414_5032.t14 a_25778_4988.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X832 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X833 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X834 a_33900_31430.t2 a_65470_24957# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.72887e+11p ps=1.96864e+06u w=1.26e+06u l=150000u
X835 a_28736_17218# a_26368_16652.t37 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X836 gnd a_56334_20860.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X837 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X838 a_26847_17217# a_23436_16644.t31 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X839 a_28736_17218# a_26368_16652.t38 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X840 a_14266_8900.t0 a_25099_11445.t40 a_17685_3840.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X841 a_23661_11500# a_14266_8900.t37 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X842 a_25815_5596# a_23414_5032.t34 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X843 a_51636_13108# Fvco_By4_QPH_bar.t8 a_51276_14152# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X844 a_28736_5597# a_26036_4988.t40 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X845 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X846 a_29252_5597# a_26036_4988.t41 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X847 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X848 vdd vdd vinit.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X849 a_45810_16322# Fvco_By4_QPH.t11 a_47760_15642# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X850 a_26073_5596# a_23414_5032.t35 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X851 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X852 a_63110_26170# a_62034_26121# a_62649_26383# gnd sky130_fd_pr__nfet_01v8 ad=2.21102e+11p pd=1.50943e+06u as=1.264e+11p ps=1.035e+06u w=640000u l=150000u
X853 a_64991_25292# a_64225_24908.t5 a_64835_25020# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.41e+10p pd=630000u as=7.63e+10p ps=923333u w=420000u l=150000u
X854 gnd gnd vbiasr.t29 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X855 a_38070_8852.t1 a_25099_11445.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X856 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X857 a_33900_31430.t4 a_65470_24957# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.84926e+11p ps=1.37203e+06u w=840000u l=150000u
X858 vdd Vso2b a_4226_12188# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X859 a_23156_5032.t3 a_14188_14050.t41 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X860 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X861 a_26110_16652# a_23436_16644.t32 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X862 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X863 vinit.t29 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X864 a_23661_11500# a_14266_8900.t38 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X865 a_27962_5597# a_26036_4988.t42 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X866 a_23661_11500# a_14266_8900.t39 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X867 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X868 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X869 a_28438_10874.t3 a_27762_11446.t33 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X870 a_26331_5596# a_23414_5032.t36 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X871 a_25557_5596# a_23414_5032.t37 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X872 a_55602_11692# Fvco_By4_QPH_bar.t9 a_50320_14126# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X873 gnd a_17685_3840.t44 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X874 a_28478_5597# a_26036_4988.t43 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X875 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X876 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X877 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X878 a_23661_11500# a_14266_8900.t40 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X879 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X880 a_23661_5596# a_14188_14050.t42 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X881 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X882 vdd Vso3b a_4226_11996# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X883 a_26073_17217# a_23436_16644.t33 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X884 a_27762_11446.t1 a_26368_16652.t39 a_28622_16652# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X885 gnd a_17685_3840.t45 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X886 a_25778_4988.t3 a_23414_5032.t38 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X887 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X888 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X889 a_8752_10532# Vso7b a_4226_11612# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X890 gnd gnd vinit.t28 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X891 a_23661_17217# a_22429_17162.t37 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X892 a_44810_16322# Fvco_By4_QPH.t12 a_47968_16078# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X893 a_62146_26505# a_62307_26207# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.155e+11p pd=1.39e+06u as=9.09625e+10p ps=656213u w=420000u l=150000u
X894 a_4314_12140# a_4288_12110# a_4314_12044# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X895 a_26331_17217# a_23436_16644.t34 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X896 a_28438_10874.t2 a_27762_11446.t34 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X897 a_56602_11692# a_51636_13108# a_52052_20860.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X898 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X899 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X900 a_25557_11500# a_25099_11445.t42 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X901 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X902 gnd a_17685_3840.t46 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X903 a_26331_17217# a_23436_16644.t35 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X904 a_28438_10874.t1 a_27762_11446.t35 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X905 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X906 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X907 vdd a_63110_26170# a_63282_26362# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=5.88e+10p ps=700000u w=420000u l=150000u
X908 a_25557_11500# a_25099_11445.t43 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X909 a_22429_17162.t0 a_26036_4988.t44 a_17685_3840.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X910 a_25299_5596# a_23414_5032.t39 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X911 a_23403_11500# a_14266_8900.t41 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X912 a_28438_10874.t0 a_27762_11446.t36 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X913 a_55602_11692# Fvco_By4_QPH_bar.t10 a_51334_14126# gnd sky130_fd_pr__nfet_01v8 ad=1.98421e+11p pd=1.49053e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X914 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X915 a_25299_11500# a_25099_11445.t44 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X916 a_26847_5596# a_23414_5032.t40 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X917 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X918 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X919 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X920 vdd vdd vinit.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X921 a_28622_16652# a_26368_16652.t40 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X922 a_25557_17217# a_23436_16644.t36 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X923 a_24177_11500# a_14266_8900.t42 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X924 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X925 a_28220_5597# a_26036_4988.t45 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X926 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X927 a_64884_26512# Fvco_By4_QPH.t13 a_65003_26240# gnd sky130_fd_pr__nfet_01v8 ad=1.134e+11p pd=960000u as=4.41e+10p ps=630000u w=420000u l=150000u
X928 a_26690_784.t1 a_23414_5032.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X929 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X930 a_29252_11501# a_27762_11446.t37 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X931 a_24177_11500# a_14266_8900.t43 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X932 a_23403_11500# a_14266_8900.t44 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X933 a_77598_24640.t3 a_77572_23336.t1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X934 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X935 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X936 gnd gnd vinit.t27 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X937 a_29252_11501# a_27762_11446.t38 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X938 a_55602_11692# a_51041_13108# a_52052_20860.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X939 a_26073_5596# a_23414_5032.t42 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X940 a_23403_11500# a_14266_8900.t45 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X941 vbiasbuffer.t1 vbiasbuffer.t0 a_54452_7044.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X942 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X943 a_65437_26240# a_65387_26390# a_65360_26240# gnd sky130_fd_pr__nfet_01v8 ad=5.775e+10p pd=695000u as=4.935e+10p ps=655000u w=420000u l=150000u
X944 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X945 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X946 a_24177_17217# a_22429_17162.t38 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X947 a_23403_11500# a_14266_8900.t46 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X948 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X949 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X950 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X951 a_25815_17217# a_23436_16644.t37 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X952 a_47760_15642# Fvco_By4_QPH_bar.t11 a_45810_16322# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.33143e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X953 a_26589_5596# a_23414_5032.t43 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X954 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X955 a_26847_17217# a_23436_16644.t38 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X956 a_14188_14050.t0 a_14266_8900.t47 a_23160_10936.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X957 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X958 gnd a_4226_12188# a_4314_12140# gnd sky130_fd_pr__nfet_01v8 ad=7.13285e+11p pd=5.29211e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X959 vdd Vso5b a_4226_11804# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X960 a_29252_17218# a_26368_16652.t41 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X961 vbiasr.t7 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X962 a_23403_17217# a_22429_17162.t39 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X963 a_26847_17217# a_23436_16644.t39 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X964 a_28478_11501# a_27762_11446.t39 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X965 a_50112_7696# a_54394_7696# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X966 a_51334_14126# Fvco_By4_QPH.t14 a_55602_11692# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X967 a_53276_4354# a_49858_3690.t9 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.856e+11p pd=1.57e+06u as=2.81792e+11p ps=2.09071e+06u w=1.28e+06u l=8e+06u
X968 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X969 gnd a_17685_3840.t47 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X970 Vso2b a_28790_25040.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X971 a_62475_26233# a_61865_26121.t5 a_62146_26505# gnd sky130_fd_pr__nfet_01v8 ad=1.2285e+11p pd=1.005e+06u as=1.134e+11p ps=960000u w=420000u l=150000u
X972 a_66020_26369# a_65848_26177# a_66158_26177# gnd sky130_fd_pr__nfet_01v8 ad=1.113e+11p pd=1.37e+06u as=4.41e+10p ps=630000u w=420000u l=150000u
X973 vinit.t26 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X974 a_29252_17218# a_26368_16652.t42 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X975 a_47760_15642# Fvco_By4_QPH_bar.t12 a_44810_16322# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X976 a_22972_23306.t4 a_23504_23306# gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X977 a_28478_11501# a_27762_11446.t40 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X978 a_50262_14152# a_50320_14126# a_50511_16072.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X979 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X980 a_23919_11500# a_14266_8900.t48 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X981 a_28478_11501# a_27762_11446.t41 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X982 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X983 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X984 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X985 a_23919_11500# a_14266_8900.t49 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X986 a_28478_11501# a_27762_11446.t42 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X987 vdd vdd vbiasr.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X988 a_26331_5596# a_23414_5032.t44 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X989 gnd gnd vbiasr.t28 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X990 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X991 a_63240_26538# a_62034_26121# a_63110_26170# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.41e+10p pd=630000u as=8.96e+10p ps=810000u w=420000u l=150000u
X992 a_23661_17217# a_22429_17162.t40 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X993 a_22887_11500# a_14266_8900.t50 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X994 a_47968_16078# Fvco_By4_QPH_bar.t13 a_45810_16322# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X995 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X996 vinit.t6 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X997 Vso1b a_24410_25128.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X998 a_28478_17218# a_26368_16652.t43 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X999 a_23661_17217# a_22429_17162.t41 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1000 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1001 a_23919_17217# a_22429_17162.t42 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1002 a_22887_11500# a_14266_8900.t51 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1003 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1004 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1005 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1006 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1007 a_62034_26121# a_61865_26121.t6 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.696e+11p pd=1.81e+06u as=1.38609e+11p ps=999944u w=640000u l=150000u
X1008 a_42550_16062# Fvco_By4_QPH.t15 a_42782_16060# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X1009 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1010 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1011 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1012 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1013 a_22887_17217# a_22429_17162.t43 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1014 vdd vdd vbiasr.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1015 Vso4b a_38070_8852.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X1016 a_52052_20860.t2 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X1017 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1018 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1019 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1020 a_28622_16652# a_26368_16652.t44 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1021 a_23145_5596# a_14188_14050.t43 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1022 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1023 gnd a_62307_26207# a_64225_24908.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=0p ps=0u w=420000u l=150000u
X1024 a_25557_17217# a_23436_16644.t40 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1025 vdd a_4288_11534# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1026 a_28622_16652# a_26368_16652.t45 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1027 a_65003_26240# reset gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=9.24629e+10p ps=686014u w=420000u l=150000u
X1028 a_17685_3840.t2 vctrl a_22972_23306.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1029 a_25557_17217# a_23436_16644.t41 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1030 gnd gnd vbiasr.t27 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1031 a_62307_26207# a_63110_26170# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.764e+11p pd=1.54e+06u as=2.72887e+11p ps=1.96864e+06u w=1.26e+06u l=150000u
X1032 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1033 vdd a_64066_26111# a_64603_26128.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38609e+11p pd=999944u as=0p ps=0u w=640000u l=150000u
X1034 a_77280_24640.t3 a_77254_23336.t2 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1035 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1036 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1037 a_23145_17217# a_22429_17162.t44 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1038 a_24177_17217# a_22429_17162.t45 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1039 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1040 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1041 gnd a_17685_3840.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1042 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1043 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1044 gnd gnd vinit.t25 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1045 a_24177_17217# a_22429_17162.t46 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1046 gnd a_17685_3840.t49 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1047 a_29252_17218# a_26368_16652.t46 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1048 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1049 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1050 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1051 a_23403_17217# a_22429_17162.t47 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1052 a_22887_5596# a_14188_14050.t44 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1053 vbiasbuffer.t2 a_49858_3690.t10 a_54950_2532# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.175e+11p ps=1.79e+06u w=1.5e+06u l=8e+06u
X1054 a_52052_20860.t11 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X1055 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1056 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1057 a_29252_17218# a_26368_16652.t47 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1058 a_23403_17217# a_22429_17162.t48 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1059 a_26589_11500# a_25099_11445.t45 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1060 a_22629_11500# a_14266_8900.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1061 a_54950_2532# a_49858_3690.t11 a_53292_2532# gnd sky130_fd_pr__nfet_01v8 ad=2.175e+11p pd=1.79e+06u as=2.175e+11p ps=1.79e+06u w=1.5e+06u l=8e+06u
X1062 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1063 a_17685_3840.t4 vinit.t40 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16577e+11p ps=1.56241e+06u w=1e+06u l=2e+06u
X1064 a_24177_5596# a_14188_14050.t45 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1065 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1066 a_22629_11500# a_14266_8900.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1067 vdd a_65387_26390# a_65369_26512# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=4.41e+10p ps=630000u w=420000u l=150000u
X1068 vdd vdd vbiasr.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1069 a_50511_16072.t6 a_42550_16062# a_47968_16078# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1070 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1071 vdd a_51138_20858# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1072 gnd a_17685_3840.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1073 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1074 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1075 a_62649_26383# a_62475_26233# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.264e+11p pd=1.035e+06u as=1.40896e+11p ps=1.04535e+06u w=640000u l=150000u
X1076 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1077 a_22629_17217# a_22429_17162.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1078 Vso6b a_14832_12082.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X1079 vdd Vso4b a_4226_11996# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1080 a_26589_11500# a_25099_11445.t46 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1081 a_28994_5597# a_26036_4988.t46 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1082 a_56602_11692# a_51636_13108# a_52052_20860.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1083 a_50511_16072.t2 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1084 a_51276_14152# Fvco_By4_QPH.t16 a_51041_13108# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1085 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1086 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1087 vinit.t5 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1088 a_26589_11500# a_25099_11445.t47 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1089 Fvco_By4_QPH_bar.t0 a_66604_26416# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.72887e+11p ps=1.96864e+06u w=1.26e+06u l=150000u
X1090 a_65470_24957# a_64394_24908# a_65009_25170# gnd sky130_fd_pr__nfet_01v8 ad=2.21102e+11p pd=1.50943e+06u as=1.264e+11p ps=1.035e+06u w=640000u l=150000u
X1091 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1092 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1093 a_26589_11500# a_25099_11445.t48 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1094 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1095 a_28478_17218# a_26368_16652.t48 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1096 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1097 gnd gnd vbiasr.t26 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1098 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1099 a_34044_31208# a_33804_31120.t8 vctrl vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X1100 vdd Vso1b a_4226_12188# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1101 a_26589_17217# a_23436_16644.t42 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1102 a_23919_17217# a_22429_17162.t50 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1103 a_28478_17218# a_26368_16652.t49 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1104 a_28994_11501# a_27762_11446.t43 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1105 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1106 Fvco_By4_QPH.t2 a_65848_26177# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.84926e+11p ps=1.37203e+06u w=840000u l=150000u
X1107 a_64982_25020# a_64394_24908# a_64835_25020# gnd sky130_fd_pr__nfet_01v8 ad=4.935e+10p pd=655000u as=1.2285e+11p ps=1.005e+06u w=420000u l=150000u
X1108 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1109 a_56602_11692# Fvco_By4_QPH_bar.t14 a_51334_14126# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1110 a_23919_17217# a_22429_17162.t51 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1111 a_43010_16058# Fvco_By4_QPH.t17 a_42782_16060# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1112 a_55602_11692# a_51041_13108# a_52052_20860.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1113 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1114 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1115 vctrl a_33900_31430.t10 a_9354_33563# vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X1116 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1117 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1118 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1119 a_24410_25128.t1 a_23436_16644.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X1120 a_22887_17217# a_22429_17162.t52 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1121 a_27962_5597# a_26036_4988.t47 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1122 vdd vdd vbiasr.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1123 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1124 a_22887_17217# a_22429_17162.t53 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1125 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1126 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1127 gnd a_17685_3840.t51 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1128 a_22629_5596# a_14188_14050.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1129 gnd a_17685_3840.t52 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1130 a_23145_5596# a_14188_14050.t47 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1131 a_23661_5596# a_14188_14050.t48 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1132 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.0821e+12p pd=2.28671e+07u as=3.0821e+12p ps=2.28671e+07u w=1.4e+07u l=1e+06u
X1133 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.2015e+11p pd=1.63337e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1134 a_45810_16322# a_77572_23336.t4 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1135 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1136 a_28790_25040.t1 a_26368_16652.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X1137 a_65642_25149# reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=9.09625e+10p ps=656213u w=420000u l=150000u
X1138 a_25299_11500# a_25099_11445.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1139 gnd a_57710_5326.t1 a_57710_5326.t2 gnd sky130_fd_pr__nfet_01v8 ad=6.60449e+11p pd=4.9001e+06u as=0p ps=0u w=3e+06u l=1e+06u
X1140 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1141 a_66020_26369# reset vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=9.09625e+10p ps=656213u w=420000u l=150000u
X1142 Vso8b a_30384_802.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.24629e+10p ps=686014u w=420000u l=150000u
X1143 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1144 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1145 a_65009_25170# a_64835_25020# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.264e+11p pd=1.035e+06u as=1.40896e+11p ps=1.04535e+06u w=640000u l=150000u
X1146 vdd Vso2b a_4288_12110# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1147 a_46856_19268.t0 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1148 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1149 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1150 vdd Vso4b a_4288_11918# vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1151 a_56602_11692# a_51636_13108# a_52052_20860.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1152 gnd a_17685_3840.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1153 a_42782_16060# a_45810_16322# a_44752_16348.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1154 vdd a_65470_24957# a_65642_25149# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=5.88e+10p ps=700000u w=420000u l=150000u
X1155 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1156 a_8748_11114# Vso6b a_4288_11726# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1157 a_26331_17217# a_23436_16644.t44 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1158 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1159 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1160 a_28736_5597# a_26036_4988.t48 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1161 a_22629_5596# a_14188_14050.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1162 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1163 a_25299_11500# a_25099_11445.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1164 vbiasr.t25 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1165 a_22887_5596# a_14188_14050.t50 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1166 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1167 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1168 vdd vdd vinit.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1169 a_62699_26233# a_62649_26383# a_62622_26233# gnd sky130_fd_pr__nfet_01v8 ad=5.775e+10p pd=695000u as=4.935e+10p ps=655000u w=420000u l=150000u
X1170 a_25299_11500# a_25099_11445.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1171 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1172 a_23919_5596# a_14188_14050.t51 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1173 a_28736_11501# a_27762_11446.t44 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1174 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1175 a_27962_11501# a_27762_11446.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1176 a_25299_11500# a_25099_11445.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1177 a_23156_5032.t2 a_14188_14050.t52 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1178 vdd reset a_64506_25292# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X1179 a_77572_23336.t6 a_77254_23336.t5 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1180 a_14188_14050.t1 a_14266_8900.t54 a_17685_3840.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1181 a_27962_11501# a_27762_11446.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1182 a_55602_11692# a_51041_13108# a_52052_20860.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1183 a_51334_14126# Fvco_By4_QPH.t18 a_56602_11692# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=1.98421e+11p ps=1.49053e+06u w=1e+06u l=150000u
X1184 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1185 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1186 a_25299_17217# a_23436_16644.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1187 a_22629_17217# a_22429_17162.t54 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1188 gnd a_17685_3840.t54 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1189 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1190 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1191 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1192 a_42574_15624# a_44810_16322# a_44752_16348.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1193 vdd a_65470_24957# a_33900_31430.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=2.72887e+11p pd=1.96864e+06u as=0p ps=0u w=1.26e+06u l=150000u
X1194 a_26073_5596# a_23414_5032.t45 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1195 a_28736_5597# a_26036_4988.t49 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1196 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1197 a_24410_25128.t0 a_23436_16644.t46 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X1198 gnd a_65470_24957# a_66226_25196# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X1199 vdd a_4288_11726# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1200 a_14832_12082.t1 a_14188_14050.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X1201 a_22629_17217# a_22429_17162.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1202 a_28478_5597# a_26036_4988.t50 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1203 a_28994_5597# a_26036_4988.t51 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1204 a_23160_10936.t2 a_14266_8900.t55 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1205 a_42574_15624# Fvco_By4_QPH_bar.t15 a_43010_16058# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1206 a_27962_17218# a_26368_16652.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1207 a_25778_4988.t2 a_23414_5032.t46 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1208 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1209 a_25099_11445.t1 a_27762_11446.t47 a_17685_3840.t9 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1210 a_23160_10936.t1 a_14266_8900.t56 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1211 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1212 a_22972_23306.t1 vctrl a_17685_3840.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1213 a_23156_5032.t1 a_14188_14050.t54 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1214 vbiasr.t24 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1215 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1216 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1217 a_17685_3840.t1 vctrl a_22972_23306.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1218 a_26589_17217# a_23436_16644.t47 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1219 vdd a_54452_7044.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1220 a_8740_12844# Vso3b a_4226_11996# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1221 a_4314_11468# a_4226_11420# v9m gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=1.0044e+12p ps=7.1e+06u w=3.24e+06u l=150000u
X1222 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1223 a_27762_11446.t0 a_26368_16652.t52 a_17685_3840.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1224 a_26589_17217# a_23436_16644.t48 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1225 a_38070_8852.t0 a_25099_11445.t53 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.19118e+11p ps=859327u w=550000u l=8e+06u
X1226 a_23178_16644# a_22429_17162.t56 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1227 a_27962_17218# a_26368_16652.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1228 a_28478_5597# a_26036_4988.t52 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1229 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1230 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1231 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1232 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1233 a_22972_23306.t3 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X1234 a_51041_13108# Fvco_By4_QPH_bar.t16 a_50262_14152# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1235 a_25778_4988.t1 a_23414_5032.t47 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1236 a_62475_26233# a_62034_26121# a_62146_26505# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.63e+10p pd=923333u as=1.155e+11p ps=1.39e+06u w=420000u l=150000u
X1237 gnd reset a_65059_25020# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=5.775e+10p ps=695000u w=420000u l=150000u
X1238 a_26847_5596# a_23414_5032.t48 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1239 a_32948_24994.t1 a_27762_11446.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=150000u
X1240 gnd a_66604_26416# Fvco_By4_QPH_bar.t2 gnd sky130_fd_pr__nfet_01v8 ad=1.84926e+11p pd=1.37203e+06u as=0p ps=0u w=840000u l=150000u
X1241 a_28578_5014.t1 a_26036_4988.t53 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1242 vbiasr.t23 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1243 a_65622_24957# a_64225_24908.t6 a_65470_24957# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.45098e+11p ps=990566u w=420000u l=150000u
X1244 a_28220_5597# a_26036_4988.t54 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1245 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1246 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1247 a_65600_25325# a_64394_24908# a_65470_24957# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.41e+10p pd=630000u as=8.96e+10p ps=810000u w=420000u l=150000u
X1248 a_22629_5596# a_14188_14050.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1249 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1250 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1251 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1252 a_55602_11692# vbiasob.t4 a_51138_21494.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=2e+06u
X1253 a_23403_5596# a_14188_14050.t56 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1254 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1255 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1256 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1257 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1258 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1259 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1260 a_63110_26170# a_61865_26121.t7 a_62649_26383# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.792e+11p pd=1.62e+06u as=2.41013e+11p ps=1.515e+06u w=840000u l=150000u
X1261 gnd a_65470_24957# a_33900_31430.t3 gnd sky130_fd_pr__nfet_01v8 ad=1.84926e+11p pd=1.37203e+06u as=0p ps=0u w=840000u l=150000u
X1262 vdd a_4226_11612# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1263 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1264 a_64394_24908# a_64225_24908.t7 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.696e+11p pd=1.81e+06u as=1.38609e+11p ps=999944u w=640000u l=150000u
X1265 a_23661_17217# a_22429_17162.t57 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1266 a_51041_13108# Fvco_By4_QPH_bar.t17 a_51276_14152# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.07143e+11p ps=1.67714e+06u w=1e+06u l=150000u
X1267 a_26847_5596# a_23414_5032.t49 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1268 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1269 a_26589_5596# a_23414_5032.t50 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1270 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1271 a_28220_5597# a_26036_4988.t55 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1272 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1273 a_4314_11852# a_4226_11804# a_4314_11756# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X1274 a_26016_10878.t1 a_25099_11445.t54 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1275 a_26016_10878.t0 a_25099_11445.t55 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1276 a_28736_5597# a_26036_4988.t56 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1277 a_29510_5597# a_26036_4988.t57 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1278 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1279 gnd a_63110_26170# a_63866_26409# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=1.113e+11p ps=1.37e+06u w=420000u l=150000u
X1280 a_44810_16322# vbiasbuffer.t4 a_50032_16080.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=1e+06u
X1281 vbiasr.t22 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1282 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1283 a_26847_11500# a_25099_11445.t56 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1284 a_51636_13108# Fvco_By4_QPH_bar.t18 a_50262_14152# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.07143e+11p ps=1.67714e+06u w=1e+06u l=150000u
X1285 a_66158_26177# reset gnd gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=9.24629e+10p ps=686014u w=420000u l=150000u
X1286 a_8748_11692# Vso5b a_4226_11804# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1287 a_26073_11500# a_25099_11445.t57 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1288 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1289 a_50262_14152# Fvco_By4_QPH.t19 a_51636_13108# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1290 a_23156_5032.t0 a_14188_14050.t57 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1291 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1292 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1293 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1294 a_8744_9386# Fvco a_4226_11420# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1295 gnd a_17685_3840.t55 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1296 a_26589_5596# a_23414_5032.t51 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1297 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1298 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1299 a_26110_16652# a_23436_16644.t49 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1300 a_25299_17217# a_23436_16644.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1301 a_26073_11500# a_25099_11445.t58 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1302 vbiasr.t21 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1303 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1304 vdd a_66226_25196# a_33804_31120.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=2.72887e+11p pd=1.96864e+06u as=0p ps=0u w=1.26e+06u l=150000u
X1305 gnd a_65642_25149# a_65622_24957# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=4.41e+10p ps=630000u w=420000u l=150000u
X1306 a_25299_17217# a_23436_16644.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1307 vbiasr.t2 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1308 gnd a_17685_3840.t56 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1309 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1310 a_44752_16348.t3 a_45810_16322# a_42782_16060# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1311 a_25815_5596# a_23414_5032.t52 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1312 vdd a_62649_26383# a_62631_26505# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=4.41e+10p ps=630000u w=420000u l=150000u
X1313 vdd a_65642_25149# a_65600_25325# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.09625e+10p pd=656213u as=4.41e+10p ps=630000u w=420000u l=150000u
X1314 a_27962_17218# a_26368_16652.t54 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1315 a_26331_5596# a_23414_5032.t53 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1316 gnd a_17685_3840.t57 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1317 a_28478_5597# a_26036_4988.t58 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1318 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1319 gnd Vso8b a_8752_10532# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1320 a_29252_5597# a_26036_4988.t59 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1321 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1322 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1323 a_26073_17217# a_23436_16644.t52 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1324 a_27962_17218# a_26368_16652.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1325 a_25778_4988.t0 a_23414_5032.t54 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1326 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1327 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1328 a_47760_15642# a_43010_16058# a_33808_31746# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.08286e+07u as=9.47286e+11p ps=7.07857e+06u w=5e+06u l=1e+06u
X1329 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1330 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1331 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1332 a_23403_17217# a_22429_17162.t58 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1333 a_4314_11948# a_4288_11918# a_4314_11852# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X1334 gnd a_17685_3840.t58 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1335 a_23178_16644# a_22429_17162.t59 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1336 a_77598_24640.t4 a_77572_23336.t0 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1337 a_23178_16644# a_22429_17162.t60 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1338 a_25557_5596# a_23414_5032.t55 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1339 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1340 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1341 a_44752_16348.t0 a_44810_16322# a_42574_15624# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1342 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1343 a_26331_5596# a_23414_5032.t56 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1344 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.416e+07u w=2.4e+07u
X1345 vinit.t24 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1346 gnd Vso6b a_8748_11692# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1347 a_28994_11501# a_27762_11446.t49 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1348 vbiasr.t1 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1349 a_26847_5596# a_23414_5032.t57 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1350 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1351 a_54934_4354# a_49858_3690.t12 a_53276_4354# gnd sky130_fd_pr__nfet_01v8 ad=1.856e+11p pd=1.57e+06u as=1.856e+11p ps=1.57e+06u w=1.28e+06u l=8e+06u
X1352 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1353 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1354 a_25815_11500# a_25099_11445.t59 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1355 a_28220_5597# a_26036_4988.t60 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1356 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1357 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1358 Fvco_By4_QPH.t0 a_65848_26177# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.72887e+11p ps=1.96864e+06u w=1.26e+06u l=150000u
X1359 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1360 vdd a_63110_26170# a_63866_26409# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38609e+11p pd=999944u as=1.696e+11p ps=1.81e+06u w=640000u l=150000u
X1361 a_25815_11500# a_25099_11445.t60 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1362 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1363 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1364 vinit.t23 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.10075e+12p ps=8.16683e+06u w=5e+06u l=1e+06u
X1365 a_8748_9956# Vso8b a_4288_11534# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1366 gnd a_17685_3840.t59 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1367 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1368 a_25557_11500# a_25099_11445.t61 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1369 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1370 a_28994_11501# a_27762_11446.t50 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1371 a_25299_5596# a_23414_5032.t58 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.2015e+11p ps=1.63337e+06u w=1e+06u l=1e+06u
X1372 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1373 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1374 vinit.t3 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1375 a_28994_11501# a_27762_11446.t51 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1376 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1377 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1378 vdd a_4288_12110# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1379 a_25815_17217# a_23436_16644.t53 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1380 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1381 a_26589_5596# a_23414_5032.t59 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1382 a_28994_11501# a_27762_11446.t52 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1383 Vso8b a_30384_802.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.6385e+11p ps=2.62485e+06u w=1.68e+06u l=150000u
X1384 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1385 a_29510_11501# a_27762_11446.t53 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1386 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1387 a_24177_11500# a_14266_8900.t57 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1388 a_33808_31746# a_43010_16058# a_47760_15642# vdd sky130_fd_pr__pfet_01v8_lvt ad=9.47286e+11p pd=7.07857e+06u as=1.45e+12p ps=1.08286e+07u w=5e+06u l=1e+06u
X1389 a_44810_16322# a_77254_23336.t6 gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1390 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1391 a_29510_11501# a_27762_11446.t54 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1392 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1393 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1394 a_28994_17218# a_26368_16652.t56 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1395 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1396 gnd a_17685_3840.t60 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.54105e+12p pd=1.14336e+07u as=1.54105e+12p ps=1.14336e+07u w=7e+06u l=8e+06u
X1397 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1398 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1399 a_65369_26512# a_64603_26128.t7 a_65213_26240# vdd sky130_fd_pr__pfet_01v8_hvt ad=4.41e+10p pd=630000u as=7.63e+10p ps=923333u w=420000u l=150000u
X1400 a_29252_11501# a_27762_11446.t55 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1401 a_42782_16060# Fvco_By4_QPH_bar.t19 a_42550_16062# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1402 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1403 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1404 a_26110_16652# a_23436_16644.t54 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1405 a_50320_14126# Fvco_By4_QPH.t20 a_56602_11692# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X1406 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1407 a_29510_17218# a_26368_16652.t57 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1408 a_62649_26383# a_62475_26233# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.41013e+11p pd=1.515e+06u as=1.81925e+11p ps=1.31243e+06u w=840000u l=150000u
X1409 a_26110_16652# a_23436_16644.t55 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1410 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1411 gnd reset a_65437_26240# gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=5.775e+10p ps=695000u w=420000u l=150000u
X1412 a_28736_11501# a_27762_11446.t56 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1413 vdd a_54394_7696# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1414 a_50262_14152# a_50320_14126# a_50511_16072.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X1415 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1416 vdd vdd vinit.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1417 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1418 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1419 a_26073_17217# a_23436_16644.t56 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1420 a_51276_14152# a_51334_14126# a_33808_31746# gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=3.78571e+11p ps=2.99714e+06u w=2e+06u l=1e+06u
X1421 a_26331_5596# a_23414_5032.t60 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1422 gnd gnd vinit.t22 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1423 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1424 a_26073_17217# a_23436_16644.t57 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1425 vdd a_4226_11804# v9m vdd sky130_fd_pr__pfet_01v8 ad=3.6385e+11p pd=2.62485e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1426 a_29510_17218# a_26368_16652.t58 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1427 vbiasob.t2 a_57710_5326.t5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.24553e+11p ps=1.66603e+06u w=1.02e+06u l=1e+06u
X1428 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1429 a_28736_11501# a_27762_11446.t57 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1430 vbiasr.t0 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1431 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1432 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1433 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1434 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1435 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1436 a_28736_11501# a_27762_11446.t58 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1437 a_23919_5596# a_14188_14050.t58 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1438 a_50511_16072.t0 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1439 gnd gnd vinit.t21 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1440 a_28736_11501# a_27762_11446.t59 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1441 a_23919_11500# a_14266_8900.t58 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1442 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1443 a_8736_14034# Vso1b a_4226_12188# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1444 vdd vdd vinit.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08289e+12p pd=7.81206e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1445 a_28736_17218# a_26368_16652.t59 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1446 a_23145_11500# a_14266_8900.t59 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1447 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1448 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1449 a_23145_5596# a_14188_14050.t59 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1450 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1451 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1452 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1453 a_23145_11500# a_14266_8900.t60 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1454 gnd gnd vbiasr.t20 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1455 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1456 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1457 gnd Fvco a_8748_9956# gnd sky130_fd_pr__nfet_01v8 ad=1.62911e+11p pd=1.20869e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1458 a_28220_11501# a_27762_11446.t60 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1459 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1460 gnd gnd vinit.t20 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.10075e+12p pd=8.16683e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1461 a_22887_11500# a_14266_8900.t61 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1462 a_28220_11501# a_27762_11446.t61 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1463 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1464 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1465 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1466 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1467 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1468 a_23145_17217# a_22429_17162.t61 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1469 a_77280_24640.t4 a_77254_23336.t1 sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1470 gnd Fvco a_61865_26121.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.24629e+10p pd=686014u as=0p ps=0u w=420000u l=150000u
X1471 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=2.363e+07u
X1472 a_25815_17217# a_23436_16644.t58 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1473 a_33808_31746# a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=3.78571e+11p pd=2.99714e+06u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1474 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1475 a_28220_17218# a_26368_16652.t60 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1476 a_26589_17217# a_23436_16644.t59 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1477 a_26368_16652.t0 a_23436_16644.t60 a_17685_3840.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1478 a_25815_17217# a_23436_16644.t61 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1479 a_23145_5596# a_14188_14050.t60 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1480 a_8744_13422# Vso2b a_4288_12110# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1481 a_22887_5596# a_14188_14050.t61 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1482 a_44810_16322# Fvco_By4_QPH.t21 a_47760_15642# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.33143e+06u w=2e+06u l=150000u
X1483 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1484 vinit.t0 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08289e+12p ps=7.81206e+06u w=5e+06u l=1e+06u
X1485 a_8748_12270# Vso4b a_4288_11918# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1486 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1487 a_28994_17218# a_26368_16652.t61 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1488 a_28578_5014.t0 a_26036_4988.t61 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1489 vdd a_34044_31208# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
X1490 vdd a_9354_33563# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51604e+12p pd=1.09369e+07u as=1.51604e+12p ps=1.09369e+07u w=7e+06u l=8e+06u
C0 a_4226_12188# v9m 2.67fF
C1 a_56602_11692# a_51334_14126# 2.10fF
C2 a_44810_16322# a_47968_16078# 3.02fF
C3 Vso1b Vso2b 3.79fF
C4 Vso7b Vso8b 12.19fF
C5 a_4288_11534# vdd 2.42fF
C6 a_55602_11692# a_56602_11692# 2.04fF
C7 Fvco Vso4b 27.27fF
C8 Vso1b vdd 3.70fF
C9 a_42574_15624# a_43010_16058# 2.25fF
C10 a_42550_16062# a_42574_15624# 2.35fF
C11 a_4226_11804# vdd 2.43fF
C12 a_51041_13108# a_51636_13108# 4.40fF
C13 vdd Vso6b 3.09fF
C14 vdd vbiasr 50.30fF
C15 Vso5b vdd 5.20fF
C16 Vso1b vctrl 3.89fF
C17 a_45810_16322# a_47760_15642# 4.36fF
C18 vinit vdd 58.74fF
C19 Fvco_By4_QPH_bar a_45810_16322# 2.30fF
C20 Vso2b vdd 3.24fF
C21 a_55602_11692# a_51334_14126# 2.35fF
C22 a_56602_11692# a_50320_14126# 2.53fF
C23 a_47760_15642# a_47968_16078# 3.20fF
C24 a_9354_33563# vdd 505.57fF
C25 a_44810_16322# a_47760_15642# 2.29fF
C26 Fvco_By4_QPH_bar Fvco_By4_QPH 14.47fF
C27 vdd a_42550_16062# 5.00fF
C28 a_4226_11420# vdd 2.26fF
C29 a_42574_15624# a_42782_16060# 2.88fF
C30 a_42550_16062# a_43010_16058# 4.58fF
C31 Fvco vbiasr 2.24fF
C32 a_4288_11726# vdd 2.30fF
C33 a_51636_13108# a_51276_14152# 2.56fF
C34 vdd vbiasob 2.61fF
C35 vdd v9m 10.85fF
C36 a_50262_14152# a_51636_13108# 2.25fF
C37 Fvco_By4_QPH_bar vdd 2.92fF
C38 reset vdd 4.47fF
C39 Fvco vdd 5.44fF
C40 Vso3b vdd 3.96fF
C41 vdd a_4288_11918# 2.56fF
C42 a_50320_14126# a_51334_14126# 2.95fF
C43 a_34044_31208# vdd 504.99fF
C44 a_55602_11692# a_50320_14126# 2.15fF
C45 Vso7b vdd 2.92fF
C46 a_42782_16060# a_43010_16058# 2.44fF
C47 a_4226_11612# vdd 2.37fF
C48 a_51636_13108# a_56602_11692# 2.40fF
C49 vbiasot vbiasbuffer 4.18fF
C50 a_42550_16062# a_42782_16060# 2.13fF
C51 a_51041_13108# a_51276_14152# 2.50fF
C52 vdd a_4288_12110# 2.60fF
C53 vdd Vso4b 3.85fF
C54 vdd a_4226_12188# 2.55fF
C55 a_50262_14152# a_51041_13108# 4.39fF
C56 a_33808_31746# a_51334_14126# 3.18fF
C57 a_9354_33563# a_33808_31746# 2.54fF
C58 a_45810_16322# a_47968_16078# 2.43fF
C59 a_44810_16322# a_45810_16322# 2.90fF
C60 vdd a_4226_11996# 2.88fF
R0 a_26368_16652.t24 a_26368_16652.t50 1273.78
R1 a_26368_16652.n3 a_26368_16652.t52 182.777
R2 a_26368_16652.n3 a_26368_16652.t0 127.728
R3 a_26368_16652.t52 a_26368_16652.t21 113.753
R4 a_26368_16652.t52 a_26368_16652.t27 113.753
R5 a_26368_16652.t52 a_26368_16652.t43 113.753
R6 a_26368_16652.t52 a_26368_16652.t59 113.753
R7 a_26368_16652.t52 a_26368_16652.t53 113.753
R8 a_26368_16652.t52 a_26368_16652.t3 113.753
R9 a_26368_16652.t52 a_26368_16652.t16 113.753
R10 a_26368_16652.t52 a_26368_16652.t32 113.753
R11 a_26368_16652.t39 a_26368_16652.t28 113.753
R12 a_26368_16652.t39 a_26368_16652.t42 113.753
R13 a_26368_16652.t39 a_26368_16652.t58 113.753
R14 a_26368_16652.t39 a_26368_16652.t12 113.753
R15 a_26368_16652.n0 a_26368_16652.t35 113.753
R16 a_26368_16652.n0 a_26368_16652.t48 113.753
R17 a_26368_16652.t39 a_26368_16652.t6 113.753
R18 a_26368_16652.t39 a_26368_16652.t61 113.753
R19 a_26368_16652.t39 a_26368_16652.t13 113.753
R20 a_26368_16652.t39 a_26368_16652.t29 113.753
R21 a_26368_16652.t39 a_26368_16652.t44 113.753
R22 a_26368_16652.n0 a_26368_16652.t22 113.753
R23 a_26368_16652.n0 a_26368_16652.t54 113.753
R24 a_26368_16652.n0 a_26368_16652.t8 113.753
R25 a_26368_16652.n0 a_26368_16652.t19 113.753
R26 a_26368_16652.t39 a_26368_16652.t37 113.753
R27 a_26368_16652.t39 a_26368_16652.t33 113.753
R28 a_26368_16652.t39 a_26368_16652.t46 113.753
R29 a_26368_16652.t39 a_26368_16652.t4 113.753
R30 a_26368_16652.t39 a_26368_16652.t17 113.753
R31 a_26368_16652.n0 a_26368_16652.t36 113.753
R32 a_26368_16652.n1 a_26368_16652.t49 113.753
R33 a_26368_16652.n1 a_26368_16652.t7 113.753
R34 a_26368_16652.t39 a_26368_16652.t2 113.753
R35 a_26368_16652.t39 a_26368_16652.t14 113.753
R36 a_26368_16652.t39 a_26368_16652.t30 113.753
R37 a_26368_16652.t39 a_26368_16652.t45 113.753
R38 a_26368_16652.n0 a_26368_16652.t23 113.753
R39 a_26368_16652.n0 a_26368_16652.t55 113.753
R40 a_26368_16652.n0 a_26368_16652.t9 113.753
R41 a_26368_16652.n2 a_26368_16652.t20 113.753
R42 a_26368_16652.n2 a_26368_16652.t38 113.753
R43 a_26368_16652.n2 a_26368_16652.t34 113.753
R44 a_26368_16652.n2 a_26368_16652.t47 113.753
R45 a_26368_16652.n2 a_26368_16652.t5 113.753
R46 a_26368_16652.n2 a_26368_16652.t18 113.753
R47 a_26368_16652.t52 a_26368_16652.t51 113.753
R48 a_26368_16652.t52 a_26368_16652.t60 113.753
R49 a_26368_16652.t52 a_26368_16652.t15 113.753
R50 a_26368_16652.t52 a_26368_16652.t31 113.753
R51 a_26368_16652.t39 a_26368_16652.t26 113.753
R52 a_26368_16652.t39 a_26368_16652.t41 113.753
R53 a_26368_16652.t39 a_26368_16652.t57 113.753
R54 a_26368_16652.t39 a_26368_16652.t11 113.753
R55 a_26368_16652.t52 a_26368_16652.t56 113.753
R56 a_26368_16652.t52 a_26368_16652.t10 113.753
R57 a_26368_16652.t52 a_26368_16652.t25 113.753
R58 a_26368_16652.t52 a_26368_16652.t40 113.753
R59 a_26368_16652.t1 a_26368_16652.n3 57.482
R60 a_26368_16652.t52 a_26368_16652.n0 5.834
R61 a_26368_16652.t39 a_26368_16652.n1 3.384
R62 a_26368_16652.t52 a_26368_16652.t24 3.018
R63 a_26368_16652.t39 a_26368_16652.n2 2.785
R64 a_26368_16652.t52 a_26368_16652.t39 2.574
R65 a_23414_5032.t2 a_23414_5032.t41 1273.78
R66 a_23414_5032.n4 a_23414_5032.t14 345.988
R67 a_23414_5032.n3 a_23414_5032.t5 113.753
R68 a_23414_5032.n3 a_23414_5032.t3 113.753
R69 a_23414_5032.n3 a_23414_5032.t15 113.753
R70 a_23414_5032.n2 a_23414_5032.t36 113.753
R71 a_23414_5032.n2 a_23414_5032.t33 113.753
R72 a_23414_5032.n2 a_23414_5032.t31 113.753
R73 a_23414_5032.n2 a_23414_5032.t30 113.753
R74 a_23414_5032.n0 a_23414_5032.t7 113.753
R75 a_23414_5032.n0 a_23414_5032.t39 113.753
R76 a_23414_5032.n0 a_23414_5032.t37 113.753
R77 a_23414_5032.n0 a_23414_5032.t34 113.753
R78 a_23414_5032.n0 a_23414_5032.t45 113.753
R79 a_23414_5032.t14 a_23414_5032.t11 113.753
R80 a_23414_5032.t14 a_23414_5032.t8 113.753
R81 a_23414_5032.t14 a_23414_5032.t6 113.753
R82 a_23414_5032.t14 a_23414_5032.t4 113.753
R83 a_23414_5032.n0 a_23414_5032.t21 113.753
R84 a_23414_5032.n0 a_23414_5032.t17 113.753
R85 a_23414_5032.n1 a_23414_5032.t35 113.753
R86 a_23414_5032.n1 a_23414_5032.t56 113.753
R87 a_23414_5032.n1 a_23414_5032.t51 113.753
R88 a_23414_5032.n1 a_23414_5032.t49 113.753
R89 a_23414_5032.n1 a_23414_5032.t47 113.753
R90 a_23414_5032.n0 a_23414_5032.t24 113.753
R91 a_23414_5032.n0 a_23414_5032.t58 113.753
R92 a_23414_5032.n0 a_23414_5032.t55 113.753
R93 a_23414_5032.n0 a_23414_5032.t52 113.753
R94 a_23414_5032.t14 a_23414_5032.t9 113.753
R95 a_23414_5032.t14 a_23414_5032.t28 113.753
R96 a_23414_5032.t14 a_23414_5032.t25 113.753
R97 a_23414_5032.t14 a_23414_5032.t23 113.753
R98 a_23414_5032.t14 a_23414_5032.t20 113.753
R99 a_23414_5032.n0 a_23414_5032.t27 113.753
R100 a_23414_5032.t14 a_23414_5032.t26 113.753
R101 a_23414_5032.t14 a_23414_5032.t42 113.753
R102 a_23414_5032.t14 a_23414_5032.t60 113.753
R103 a_23414_5032.t14 a_23414_5032.t59 113.753
R104 a_23414_5032.t14 a_23414_5032.t57 113.753
R105 a_23414_5032.t14 a_23414_5032.t54 113.753
R106 a_23414_5032.n0 a_23414_5032.t29 113.753
R107 a_23414_5032.n0 a_23414_5032.t13 113.753
R108 a_23414_5032.n0 a_23414_5032.t12 113.753
R109 a_23414_5032.t14 a_23414_5032.t10 113.753
R110 a_23414_5032.t14 a_23414_5032.t19 113.753
R111 a_23414_5032.t14 a_23414_5032.t44 113.753
R112 a_23414_5032.t14 a_23414_5032.t43 113.753
R113 a_23414_5032.t14 a_23414_5032.t40 113.753
R114 a_23414_5032.t14 a_23414_5032.t38 113.753
R115 a_23414_5032.n0 a_23414_5032.t22 113.753
R116 a_23414_5032.n0 a_23414_5032.t18 113.753
R117 a_23414_5032.n0 a_23414_5032.t16 113.753
R118 a_23414_5032.t14 a_23414_5032.t32 113.753
R119 a_23414_5032.t14 a_23414_5032.t53 113.753
R120 a_23414_5032.t14 a_23414_5032.t50 113.753
R121 a_23414_5032.t14 a_23414_5032.t48 113.753
R122 a_23414_5032.t14 a_23414_5032.t46 113.753
R123 a_23414_5032.t0 a_23414_5032.n5 82.513
R124 a_23414_5032.n4 a_23414_5032.t1 28.697
R125 a_23414_5032.t14 a_23414_5032.n0 4.31
R126 a_23414_5032.n5 a_23414_5032.n4 3.507
R127 a_23414_5032.n0 a_23414_5032.n3 3.224
R128 a_23414_5032.t14 a_23414_5032.n1 2.869
R129 a_23414_5032.t14 a_23414_5032.n2 2.708
R130 a_23414_5032.n5 a_23414_5032.t2 2.634
R131 a_26690_784.n1 a_26690_784.t2 434.481
R132 a_26690_784.n0 a_26690_784.t3 217.163
R133 a_26690_784.t0 a_26690_784.n1 52.152
R134 a_26690_784.n0 a_26690_784.t1 3.106
R135 a_26690_784.n1 a_26690_784.n0 0.879
R136 vbiasr.n16 vbiasr.t40 11.002
R137 vbiasr.n27 vbiasr.t11 7.425
R138 vbiasr.n16 vbiasr.t10 7.425
R139 vbiasr.n25 vbiasr.t6 5.713
R140 vbiasr.n25 vbiasr.t1 5.713
R141 vbiasr.n8 vbiasr.t13 5.713
R142 vbiasr.n8 vbiasr.t2 5.713
R143 vbiasr.n9 vbiasr.t14 5.713
R144 vbiasr.n9 vbiasr.t8 5.713
R145 vbiasr.n10 vbiasr.t18 5.713
R146 vbiasr.n10 vbiasr.t9 5.713
R147 vbiasr.n11 vbiasr.t3 5.713
R148 vbiasr.n11 vbiasr.t16 5.713
R149 vbiasr.n12 vbiasr.t5 5.713
R150 vbiasr.n12 vbiasr.t17 5.713
R151 vbiasr.n13 vbiasr.t12 5.713
R152 vbiasr.n13 vbiasr.t7 5.713
R153 vbiasr.n15 vbiasr.t4 5.713
R154 vbiasr.n15 vbiasr.t0 5.713
R155 vbiasr.n14 vbiasr.t19 5.713
R156 vbiasr.n14 vbiasr.t15 5.713
R157 vbiasr.n39 vbiasr.t38 5.244
R158 vbiasr.n28 vbiasr.t37 5.244
R159 vbiasr.n0 vbiasr.t29 3.48
R160 vbiasr.n0 vbiasr.t24 3.48
R161 vbiasr.n1 vbiasr.t39 3.48
R162 vbiasr.n1 vbiasr.t25 3.48
R163 vbiasr.n2 vbiasr.t20 3.48
R164 vbiasr.n2 vbiasr.t31 3.48
R165 vbiasr.n3 vbiasr.t27 3.48
R166 vbiasr.n3 vbiasr.t35 3.48
R167 vbiasr.n4 vbiasr.t28 3.48
R168 vbiasr.n4 vbiasr.t22 3.48
R169 vbiasr.n5 vbiasr.t33 3.48
R170 vbiasr.n5 vbiasr.t23 3.48
R171 vbiasr.n6 vbiasr.t34 3.48
R172 vbiasr.n6 vbiasr.t30 3.48
R173 vbiasr.n7 vbiasr.t26 3.48
R174 vbiasr.n7 vbiasr.t36 3.48
R175 vbiasr.n29 vbiasr.t32 3.48
R176 vbiasr.n29 vbiasr.t21 3.48
R177 vbiasr.n35 vbiasr.n3 1.766
R178 vbiasr.n38 vbiasr.n0 1.766
R179 vbiasr.n32 vbiasr.n6 1.766
R180 vbiasr.n31 vbiasr.n7 1.764
R181 vbiasr.n34 vbiasr.n4 1.762
R182 vbiasr.n36 vbiasr.n2 1.761
R183 vbiasr.n33 vbiasr.n5 1.758
R184 vbiasr.n37 vbiasr.n1 1.758
R185 vbiasr.n30 vbiasr.n29 1.754
R186 vbiasr.n20 vbiasr.n12 1.714
R187 vbiasr.n17 vbiasr.n15 1.714
R188 vbiasr.n23 vbiasr.n9 1.714
R189 vbiasr.n24 vbiasr.n8 1.712
R190 vbiasr.n21 vbiasr.n11 1.71
R191 vbiasr.n19 vbiasr.n13 1.709
R192 vbiasr.n22 vbiasr.n10 1.706
R193 vbiasr.n18 vbiasr.n14 1.706
R194 vbiasr.n26 vbiasr.n25 1.702
R195 vbiasr.n28 vbiasr.n27 0.292
R196 vbiasr vbiasr.n39 0.152
R197 vbiasr.n22 vbiasr.n21 0.031
R198 vbiasr.n34 vbiasr.n33 0.031
R199 vbiasr.n19 vbiasr.n18 0.031
R200 vbiasr.n37 vbiasr.n36 0.031
R201 vbiasr.n31 vbiasr.n30 0.031
R202 vbiasr.n26 vbiasr.n24 0.031
R203 vbiasr.n30 vbiasr.n28 0.031
R204 vbiasr.n27 vbiasr.n26 0.031
R205 vbiasr.n38 vbiasr.n37 0.03
R206 vbiasr.n18 vbiasr.n17 0.03
R207 vbiasr.n39 vbiasr.n38 0.03
R208 vbiasr.n17 vbiasr.n16 0.03
R209 vbiasr.n24 vbiasr.n23 0.03
R210 vbiasr.n32 vbiasr.n31 0.03
R211 vbiasr.n21 vbiasr.n20 0.03
R212 vbiasr.n35 vbiasr.n34 0.03
R213 vbiasr.n20 vbiasr.n19 0.03
R214 vbiasr.n36 vbiasr.n35 0.03
R215 vbiasr.n33 vbiasr.n32 0.03
R216 vbiasr.n23 vbiasr.n22 0.03
R217 vinit.n18 vinit.t40 32.903
R218 vinit.n28 vinit.t12 7.425
R219 vinit.n18 vinit.t8 7.425
R220 vinit.n10 vinit.t2 5.713
R221 vinit.n10 vinit.t5 5.713
R222 vinit.n11 vinit.t10 5.713
R223 vinit.n11 vinit.t17 5.713
R224 vinit.n12 vinit.t13 5.713
R225 vinit.n12 vinit.t0 5.713
R226 vinit.n13 vinit.t4 5.713
R227 vinit.n13 vinit.t9 5.713
R228 vinit.n14 vinit.t16 5.713
R229 vinit.n14 vinit.t3 5.713
R230 vinit.n15 vinit.t7 5.713
R231 vinit.n15 vinit.t11 5.713
R232 vinit.n16 vinit.t15 5.713
R233 vinit.n16 vinit.t14 5.713
R234 vinit.n17 vinit.t1 5.713
R235 vinit.n17 vinit.t6 5.713
R236 vinit.n9 vinit.t19 5.713
R237 vinit.n9 vinit.t18 5.713
R238 vinit.n39 vinit.t24 5.244
R239 vinit.n29 vinit.t20 5.244
R240 vinit.n0 vinit.t28 3.48
R241 vinit.n0 vinit.t36 3.48
R242 vinit.n1 vinit.t35 3.48
R243 vinit.n1 vinit.t23 3.48
R244 vinit.n2 vinit.t22 3.48
R245 vinit.n2 vinit.t26 3.48
R246 vinit.n3 vinit.t34 3.48
R247 vinit.n3 vinit.t30 3.48
R248 vinit.n4 vinit.t21 3.48
R249 vinit.n4 vinit.t39 3.48
R250 vinit.n5 vinit.t25 3.48
R251 vinit.n5 vinit.t33 3.48
R252 vinit.n6 vinit.t38 3.48
R253 vinit.n6 vinit.t29 3.48
R254 vinit.n7 vinit.t27 3.48
R255 vinit.n7 vinit.t32 3.48
R256 vinit.n8 vinit.t31 3.48
R257 vinit.n8 vinit.t37 3.48
R258 vinit.n35 vinit.n3 1.766
R259 vinit.n38 vinit.n0 1.766
R260 vinit.n32 vinit.n6 1.766
R261 vinit.n31 vinit.n7 1.764
R262 vinit.n34 vinit.n4 1.762
R263 vinit.n36 vinit.n2 1.761
R264 vinit.n33 vinit.n5 1.758
R265 vinit.n37 vinit.n1 1.758
R266 vinit.n30 vinit.n8 1.754
R267 vinit.n22 vinit.n14 1.714
R268 vinit.n19 vinit.n17 1.714
R269 vinit.n25 vinit.n11 1.714
R270 vinit.n26 vinit.n10 1.712
R271 vinit.n23 vinit.n13 1.71
R272 vinit.n21 vinit.n15 1.709
R273 vinit.n24 vinit.n12 1.706
R274 vinit.n20 vinit.n16 1.706
R275 vinit.n27 vinit.n9 1.702
R276 vinit.n29 vinit.n28 0.292
R277 vinit vinit.n39 0.112
R278 vinit.n24 vinit.n23 0.031
R279 vinit.n34 vinit.n33 0.031
R280 vinit.n37 vinit.n36 0.031
R281 vinit.n21 vinit.n20 0.031
R282 vinit.n31 vinit.n30 0.031
R283 vinit.n27 vinit.n26 0.031
R284 vinit.n30 vinit.n29 0.031
R285 vinit.n28 vinit.n27 0.031
R286 vinit.n38 vinit.n37 0.03
R287 vinit.n20 vinit.n19 0.03
R288 vinit.n39 vinit.n38 0.03
R289 vinit.n19 vinit.n18 0.03
R290 vinit.n26 vinit.n25 0.03
R291 vinit.n32 vinit.n31 0.03
R292 vinit.n35 vinit.n34 0.03
R293 vinit.n23 vinit.n22 0.03
R294 vinit.n36 vinit.n35 0.03
R295 vinit.n22 vinit.n21 0.03
R296 vinit.n33 vinit.n32 0.03
R297 vinit.n25 vinit.n24 0.03
R298 a_14188_14050.t12 a_14188_14050.t53 1273.78
R299 a_14188_14050.n3 a_14188_14050.t31 161.992
R300 a_14188_14050.t39 a_14188_14050.t40 113.753
R301 a_14188_14050.t39 a_14188_14050.t50 113.753
R302 a_14188_14050.t39 a_14188_14050.t47 113.753
R303 a_14188_14050.t39 a_14188_14050.t11 113.753
R304 a_14188_14050.n0 a_14188_14050.t23 113.753
R305 a_14188_14050.n0 a_14188_14050.t6 113.753
R306 a_14188_14050.n0 a_14188_14050.t19 113.753
R307 a_14188_14050.n0 a_14188_14050.t41 113.753
R308 a_14188_14050.t39 a_14188_14050.t55 113.753
R309 a_14188_14050.t39 a_14188_14050.t9 113.753
R310 a_14188_14050.t39 a_14188_14050.t8 113.753
R311 a_14188_14050.t39 a_14188_14050.t26 113.753
R312 a_14188_14050.n0 a_14188_14050.t42 113.753
R313 a_14188_14050.n0 a_14188_14050.t24 113.753
R314 a_14188_14050.n0 a_14188_14050.t38 113.753
R315 a_14188_14050.n0 a_14188_14050.t57 113.753
R316 a_14188_14050.t31 a_14188_14050.t21 113.753
R317 a_14188_14050.t31 a_14188_14050.t36 113.753
R318 a_14188_14050.t31 a_14188_14050.t33 113.753
R319 a_14188_14050.t31 a_14188_14050.t56 113.753
R320 a_14188_14050.n0 a_14188_14050.t10 113.753
R321 a_14188_14050.n0 a_14188_14050.t51 113.753
R322 a_14188_14050.n0 a_14188_14050.t5 113.753
R323 a_14188_14050.n0 a_14188_14050.t25 113.753
R324 a_14188_14050.t31 a_14188_14050.t49 113.753
R325 a_14188_14050.t31 a_14188_14050.t4 113.753
R326 a_14188_14050.t31 a_14188_14050.t60 113.753
R327 a_14188_14050.t31 a_14188_14050.t22 113.753
R328 a_14188_14050.n1 a_14188_14050.t37 113.753
R329 a_14188_14050.n1 a_14188_14050.t18 113.753
R330 a_14188_14050.n1 a_14188_14050.t30 113.753
R331 a_14188_14050.n1 a_14188_14050.t54 113.753
R332 a_14188_14050.n2 a_14188_14050.t3 113.753
R333 a_14188_14050.n2 a_14188_14050.t16 113.753
R334 a_14188_14050.n2 a_14188_14050.t14 113.753
R335 a_14188_14050.n2 a_14188_14050.t35 113.753
R336 a_14188_14050.n0 a_14188_14050.t48 113.753
R337 a_14188_14050.n0 a_14188_14050.t29 113.753
R338 a_14188_14050.n0 a_14188_14050.t45 113.753
R339 a_14188_14050.n0 a_14188_14050.t7 113.753
R340 a_14188_14050.t31 a_14188_14050.t46 113.753
R341 a_14188_14050.t31 a_14188_14050.t61 113.753
R342 a_14188_14050.t31 a_14188_14050.t59 113.753
R343 a_14188_14050.t31 a_14188_14050.t20 113.753
R344 a_14188_14050.t31 a_14188_14050.t28 113.753
R345 a_14188_14050.t31 a_14188_14050.t44 113.753
R346 a_14188_14050.t31 a_14188_14050.t43 113.753
R347 a_14188_14050.t31 a_14188_14050.t2 113.753
R348 a_14188_14050.n0 a_14188_14050.t15 113.753
R349 a_14188_14050.n0 a_14188_14050.t58 113.753
R350 a_14188_14050.n0 a_14188_14050.t13 113.753
R351 a_14188_14050.n0 a_14188_14050.t32 113.753
R352 a_14188_14050.t31 a_14188_14050.t34 113.753
R353 a_14188_14050.t31 a_14188_14050.t17 113.753
R354 a_14188_14050.t31 a_14188_14050.t27 113.753
R355 a_14188_14050.n0 a_14188_14050.t52 113.753
R356 a_14188_14050.t0 a_14188_14050.n4 57.821
R357 a_14188_14050.n3 a_14188_14050.t1 47.07
R358 a_14188_14050.n4 a_14188_14050.t12 6.878
R359 a_14188_14050.n4 a_14188_14050.n3 3.96
R360 a_14188_14050.t31 a_14188_14050.t39 3.88
R361 a_14188_14050.t31 a_14188_14050.n0 3.25
R362 a_14188_14050.n0 a_14188_14050.n1 2.856
R363 a_14188_14050.t31 a_14188_14050.n2 2.454
R364 Fvco_By4_QPH.t12 Fvco_By4_QPH.t21 731.89
R365 Fvco_By4_QPH.t17 Fvco_By4_QPH.t9 731.89
R366 Fvco_By4_QPH.t5 Fvco_By4_QPH.t16 731.89
R367 Fvco_By4_QPH.t8 Fvco_By4_QPH.t19 718.506
R368 Fvco_By4_QPH.t14 Fvco_By4_QPH.t18 710.965
R369 Fvco_By4_QPH.t10 Fvco_By4_QPH.t17 622.637
R370 Fvco_By4_QPH.n12 Fvco_By4_QPH.n11 617.524
R371 Fvco_By4_QPH.n8 Fvco_By4_QPH.n7 580.872
R372 Fvco_By4_QPH.t18 Fvco_By4_QPH.t4 579.889
R373 Fvco_By4_QPH.n7 Fvco_By4_QPH.t15 491.229
R374 Fvco_By4_QPH.n8 Fvco_By4_QPH.t7 489.182
R375 Fvco_By4_QPH.n13 Fvco_By4_QPH.t14 418.965
R376 Fvco_By4_QPH.n12 Fvco_By4_QPH.t20 414.13
R377 Fvco_By4_QPH.n9 Fvco_By4_QPH.t11 349.273
R378 Fvco_By4_QPH.n10 Fvco_By4_QPH.t5 317.894
R379 Fvco_By4_QPH.n10 Fvco_By4_QPH.t8 291.323
R380 Fvco_By4_QPH.n9 Fvco_By4_QPH.t12 252.624
R381 Fvco_By4_QPH.n7 Fvco_By4_QPH.t10 227.612
R382 Fvco_By4_QPH.t11 Fvco_By4_QPH.n8 227.612
R383 Fvco_By4_QPH.n11 Fvco_By4_QPH.n9 198.896
R384 Fvco_By4_QPH.n13 Fvco_By4_QPH.n12 152.778
R385 Fvco_By4_QPH.n1 Fvco_By4_QPH.t6 152.326
R386 Fvco_By4_QPH.n1 Fvco_By4_QPH.t13 135.623
R387 Fvco_By4_QPH.n4 Fvco_By4_QPH.n2 42.381
R388 Fvco_By4_QPH Fvco_By4_QPH.n13 38.508
R389 Fvco_By4_QPH.n11 Fvco_By4_QPH.n10 31.687
R390 Fvco_By4_QPH.n2 Fvco_By4_QPH.t1 21.888
R391 Fvco_By4_QPH.n2 Fvco_By4_QPH.t0 21.888
R392 Fvco_By4_QPH.n3 Fvco_By4_QPH.t3 20
R393 Fvco_By4_QPH.n3 Fvco_By4_QPH.t2 20
R394 Fvco_By4_QPH Fvco_By4_QPH.n0 11.153
R395 Fvco_By4_QPH.n0 Fvco_By4_QPH.n1 9.672
R396 Fvco_By4_QPH.n4 Fvco_By4_QPH.n3 6.311
R397 Fvco_By4_QPH.n0 Fvco_By4_QPH.n6 3.988
R398 Fvco_By4_QPH.n5 Fvco_By4_QPH.n4 1.801
R399 Fvco_By4_QPH.n0 Fvco_By4_QPH.n5 0.471
R400 a_64225_24908.t3 a_64225_24908.t6 2276.65
R401 a_64225_24908.n0 a_64225_24908.t2 1000.95
R402 a_64225_24908.t7 a_64225_24908.n1 779.232
R403 a_64225_24908.n1 a_64225_24908.t4 589.347
R404 a_64225_24908.n2 a_64225_24908.t7 560.159
R405 a_64225_24908.n1 a_64225_24908.n0 298.84
R406 a_64225_24908.n0 a_64225_24908.t5 176.733
R407 a_64225_24908.t0 a_64225_24908.n3 135.884
R408 a_64225_24908.n2 a_64225_24908.t3 124.034
R409 a_64225_24908.n3 a_64225_24908.t1 62.096
R410 a_64225_24908.n3 a_64225_24908.n2 33.009
R411 a_33900_31430.n1 a_33900_31430.t10 449.587
R412 a_33900_31430.n1 a_33900_31430.t6 402.739
R413 a_33900_31430.n0 a_33900_31430.t8 270.989
R414 a_33900_31430.n0 a_33900_31430.t9 227.612
R415 a_33900_31430.n2 a_33900_31430.n0 199.119
R416 a_33900_31430.n3 a_33900_31430.t5 152.326
R417 a_33900_31430.n16 a_33900_31430.n2 138.854
R418 a_33900_31430.n3 a_33900_31430.t7 135.623
R419 a_33900_31430.t0 a_33900_31430.n16 94.674
R420 a_33900_31430.n2 a_33900_31430.n1 38.57
R421 a_33900_31430.n13 a_33900_31430.t3 20
R422 a_33900_31430.n13 a_33900_31430.t4 20
R423 a_33900_31430.n14 a_33900_31430.n13 19.705
R424 a_33900_31430.n4 a_33900_31430.t1 19.543
R425 a_33900_31430.n7 a_33900_31430.t2 10.944
R426 a_33900_31430.n15 a_33900_31430.n3 9.015
R427 a_33900_31430.n9 a_33900_31430.n8 5.496
R428 a_33900_31430.n12 a_33900_31430.n11 4.857
R429 a_33900_31430.n8 a_33900_31430.n7 4.01
R430 a_33900_31430.n8 a_33900_31430.n6 4.01
R431 a_33900_31430.n16 a_33900_31430.n15 2.761
R432 a_33900_31430.n5 a_33900_31430.n4 2.105
R433 a_33900_31430.n12 a_33900_31430.n9 0.227
R434 a_33900_31430.n6 a_33900_31430.n5 0.208
R435 a_33900_31430.n11 a_33900_31430.n10 0.139
R436 a_33900_31430.n15 a_33900_31430.n14 0.031
R437 a_33900_31430.n14 a_33900_31430.n12 0.002
R438 a_26036_4988.t16 a_26036_4988.t22 1273.78
R439 a_26036_4988.n0 a_26036_4988.t44 415.476
R440 a_26036_4988.t44 a_26036_4988.t37 113.753
R441 a_26036_4988.t44 a_26036_4988.t34 113.753
R442 a_26036_4988.t44 a_26036_4988.t32 113.753
R443 a_26036_4988.t20 a_26036_4988.t46 113.753
R444 a_26036_4988.t20 a_26036_4988.t7 113.753
R445 a_26036_4988.t20 a_26036_4988.t4 113.753
R446 a_26036_4988.t20 a_26036_4988.t61 113.753
R447 a_26036_4988.t44 a_26036_4988.t14 113.753
R448 a_26036_4988.t44 a_26036_4988.t47 113.753
R449 a_26036_4988.t44 a_26036_4988.t10 113.753
R450 a_26036_4988.t44 a_26036_4988.t6 113.753
R451 a_26036_4988.t44 a_26036_4988.t3 113.753
R452 a_26036_4988.t20 a_26036_4988.t15 113.753
R453 a_26036_4988.t20 a_26036_4988.t41 113.753
R454 a_26036_4988.t20 a_26036_4988.t38 113.753
R455 a_26036_4988.t20 a_26036_4988.t35 113.753
R456 a_26036_4988.n1 a_26036_4988.t55 113.753
R457 a_26036_4988.n1 a_26036_4988.t52 113.753
R458 a_26036_4988.t20 a_26036_4988.t49 113.753
R459 a_26036_4988.t20 a_26036_4988.t5 113.753
R460 a_26036_4988.t20 a_26036_4988.t27 113.753
R461 a_26036_4988.t20 a_26036_4988.t25 113.753
R462 a_26036_4988.t20 a_26036_4988.t18 113.753
R463 a_26036_4988.n1 a_26036_4988.t36 113.753
R464 a_26036_4988.n1 a_26036_4988.t8 113.753
R465 a_26036_4988.n1 a_26036_4988.t29 113.753
R466 a_26036_4988.n1 a_26036_4988.t26 113.753
R467 a_26036_4988.t20 a_26036_4988.t23 113.753
R468 a_26036_4988.t20 a_26036_4988.t39 113.753
R469 a_26036_4988.t20 a_26036_4988.t59 113.753
R470 a_26036_4988.t20 a_26036_4988.t57 113.753
R471 a_26036_4988.t20 a_26036_4988.t53 113.753
R472 a_26036_4988.n1 a_26036_4988.t60 113.753
R473 a_26036_4988.t20 a_26036_4988.t58 113.753
R474 a_26036_4988.t20 a_26036_4988.t56 113.753
R475 a_26036_4988.t20 a_26036_4988.t11 113.753
R476 a_26036_4988.t20 a_26036_4988.t31 113.753
R477 a_26036_4988.t20 a_26036_4988.t30 113.753
R478 a_26036_4988.t20 a_26036_4988.t28 113.753
R479 a_26036_4988.n1 a_26036_4988.t42 113.753
R480 a_26036_4988.n1 a_26036_4988.t19 113.753
R481 a_26036_4988.n1 a_26036_4988.t45 113.753
R482 a_26036_4988.n2 a_26036_4988.t43 113.753
R483 a_26036_4988.n2 a_26036_4988.t40 113.753
R484 a_26036_4988.n2 a_26036_4988.t51 113.753
R485 a_26036_4988.n2 a_26036_4988.t13 113.753
R486 a_26036_4988.n2 a_26036_4988.t12 113.753
R487 a_26036_4988.n2 a_26036_4988.t9 113.753
R488 a_26036_4988.t44 a_26036_4988.t33 113.753
R489 a_26036_4988.t44 a_26036_4988.t54 113.753
R490 a_26036_4988.t44 a_26036_4988.t50 113.753
R491 a_26036_4988.t44 a_26036_4988.t48 113.753
R492 a_26036_4988.t44 a_26036_4988.t2 113.753
R493 a_26036_4988.t44 a_26036_4988.t24 113.753
R494 a_26036_4988.t44 a_26036_4988.t21 113.753
R495 a_26036_4988.t44 a_26036_4988.t17 113.753
R496 a_26036_4988.t1 a_26036_4988.n0 81.094
R497 a_26036_4988.n0 a_26036_4988.t0 28.577
R498 a_26036_4988.t44 a_26036_4988.n1 6.49
R499 a_26036_4988.n0 a_26036_4988.t16 5.37
R500 a_26036_4988.t20 a_26036_4988.n2 4.699
R501 a_26036_4988.t44 a_26036_4988.t20 2.967
R502 a_33804_31120.n0 a_33804_31120.t8 440.519
R503 a_33804_31120.n0 a_33804_31120.t7 402.739
R504 a_33804_31120.n2 a_33804_31120.t6 227.612
R505 a_33804_31120.n1 a_33804_31120.t5 227.612
R506 a_33804_31120.n1 a_33804_31120.n0 183.872
R507 a_33804_31120.n6 a_33804_31120.n2 178.766
R508 a_33804_31120.n2 a_33804_31120.n1 45.046
R509 a_33804_31120.n5 a_33804_31120.n3 25.007
R510 a_33804_31120.n5 a_33804_31120.n4 24.147
R511 a_33804_31120.n4 a_33804_31120.t0 21.888
R512 a_33804_31120.n4 a_33804_31120.t1 21.888
R513 a_33804_31120.n3 a_33804_31120.t2 20
R514 a_33804_31120.n3 a_33804_31120.t3 20
R515 a_33804_31120.t4 a_33804_31120.n6 9.537
R516 a_33804_31120.n6 a_33804_31120.n5 3.669
R517 a_61865_26121.t4 a_61865_26121.t2 2276.65
R518 a_61865_26121.n0 a_61865_26121.t7 1000.95
R519 a_61865_26121.t6 a_61865_26121.n1 779.232
R520 a_61865_26121.n1 a_61865_26121.t5 589.347
R521 a_61865_26121.n2 a_61865_26121.t6 560.159
R522 a_61865_26121.n1 a_61865_26121.n0 298.84
R523 a_61865_26121.n0 a_61865_26121.t3 176.733
R524 a_61865_26121.t0 a_61865_26121.n3 135.884
R525 a_61865_26121.n2 a_61865_26121.t4 124.034
R526 a_61865_26121.n3 a_61865_26121.t1 62.096
R527 a_61865_26121.n3 a_61865_26121.n2 33.009
R528 a_25099_11445.t53 a_25099_11445.t41 1273.78
R529 a_25099_11445.n3 a_25099_11445.t40 218.051
R530 a_25099_11445.t40 a_25099_11445.t49 113.753
R531 a_25099_11445.t40 a_25099_11445.t8 113.753
R532 a_25099_11445.t40 a_25099_11445.t29 113.753
R533 a_25099_11445.t40 a_25099_11445.t21 113.753
R534 a_25099_11445.t40 a_25099_11445.t42 113.753
R535 a_25099_11445.t40 a_25099_11445.t59 113.753
R536 a_25099_11445.t40 a_25099_11445.t57 113.753
R537 a_25099_11445.n2 a_25099_11445.t6 113.753
R538 a_25099_11445.n2 a_25099_11445.t16 113.753
R539 a_25099_11445.n2 a_25099_11445.t37 113.753
R540 a_25099_11445.n2 a_25099_11445.t54 113.753
R541 a_25099_11445.t40 a_25099_11445.t19 113.753
R542 a_25099_11445.n0 a_25099_11445.t51 113.753
R543 a_25099_11445.n0 a_25099_11445.t10 113.753
R544 a_25099_11445.n0 a_25099_11445.t31 113.753
R545 a_25099_11445.n1 a_25099_11445.t26 113.753
R546 a_25099_11445.n1 a_25099_11445.t35 113.753
R547 a_25099_11445.n1 a_25099_11445.t47 113.753
R548 a_25099_11445.n1 a_25099_11445.t4 113.753
R549 a_25099_11445.n1 a_25099_11445.t23 113.753
R550 a_25099_11445.n0 a_25099_11445.t43 113.753
R551 a_25099_11445.n0 a_25099_11445.t60 113.753
R552 a_25099_11445.t15 a_25099_11445.t58 113.753
R553 a_25099_11445.t15 a_25099_11445.t7 113.753
R554 a_25099_11445.t15 a_25099_11445.t17 113.753
R555 a_25099_11445.t15 a_25099_11445.t38 113.753
R556 a_25099_11445.t15 a_25099_11445.t55 113.753
R557 a_25099_11445.n0 a_25099_11445.t20 113.753
R558 a_25099_11445.n0 a_25099_11445.t52 113.753
R559 a_25099_11445.n0 a_25099_11445.t11 113.753
R560 a_25099_11445.t15 a_25099_11445.t32 113.753
R561 a_25099_11445.t15 a_25099_11445.t27 113.753
R562 a_25099_11445.t15 a_25099_11445.t36 113.753
R563 a_25099_11445.t15 a_25099_11445.t48 113.753
R564 a_25099_11445.t15 a_25099_11445.t5 113.753
R565 a_25099_11445.t15 a_25099_11445.t24 113.753
R566 a_25099_11445.t15 a_25099_11445.t39 113.753
R567 a_25099_11445.t15 a_25099_11445.t56 113.753
R568 a_25099_11445.t15 a_25099_11445.t12 113.753
R569 a_25099_11445.n0 a_25099_11445.t44 113.753
R570 a_25099_11445.n0 a_25099_11445.t61 113.753
R571 a_25099_11445.t15 a_25099_11445.t14 113.753
R572 a_25099_11445.t15 a_25099_11445.t13 113.753
R573 a_25099_11445.t15 a_25099_11445.t28 113.753
R574 a_25099_11445.t40 a_25099_11445.t50 113.753
R575 a_25099_11445.t40 a_25099_11445.t9 113.753
R576 a_25099_11445.t40 a_25099_11445.t30 113.753
R577 a_25099_11445.t40 a_25099_11445.t25 113.753
R578 a_25099_11445.t15 a_25099_11445.t34 113.753
R579 a_25099_11445.t15 a_25099_11445.t46 113.753
R580 a_25099_11445.t15 a_25099_11445.t3 113.753
R581 a_25099_11445.t15 a_25099_11445.t22 113.753
R582 a_25099_11445.t40 a_25099_11445.t33 113.753
R583 a_25099_11445.t40 a_25099_11445.t45 113.753
R584 a_25099_11445.t40 a_25099_11445.t2 113.753
R585 a_25099_11445.t40 a_25099_11445.t18 113.753
R586 a_25099_11445.t0 a_25099_11445.n4 56.779
R587 a_25099_11445.n3 a_25099_11445.t1 28.581
R588 a_25099_11445.t40 a_25099_11445.n0 5.834
R589 a_25099_11445.n4 a_25099_11445.t53 4.799
R590 a_25099_11445.n4 a_25099_11445.n3 3.709
R591 a_25099_11445.t15 a_25099_11445.n1 2.869
R592 a_25099_11445.t40 a_25099_11445.t15 2.816
R593 a_25099_11445.t15 a_25099_11445.n2 2.586
R594 a_17685_3840.n27 a_17685_3840.n26 660.793
R595 a_17685_3840.n55 a_17685_3840.n54 649.743
R596 a_17685_3840.n60 a_17685_3840.n59 574.593
R597 a_17685_3840.n28 a_17685_3840.n27 416.406
R598 a_17685_3840.n61 a_17685_3840.n60 415.789
R599 a_17685_3840.n57 a_17685_3840.n56 271.45
R600 a_17685_3840.n59 a_17685_3840.n58 262.496
R601 a_17685_3840.n27 a_17685_3840.n25 198.935
R602 a_17685_3840.n59 a_17685_3840.t0 197.212
R603 a_17685_3840.n58 a_17685_3840.t7 185.816
R604 a_17685_3840.n26 a_17685_3840.t12 176.327
R605 a_17685_3840.n57 a_17685_3840.t6 173.989
R606 a_17685_3840.n25 a_17685_3840.t9 154.605
R607 a_17685_3840.n56 a_17685_3840.t8 151.674
R608 a_17685_3840.n62 a_17685_3840.t11 118.032
R609 a_17685_3840.n60 a_17685_3840.n57 107.97
R610 a_17685_3840.n29 a_17685_3840.n28 104.297
R611 a_17685_3840.n63 a_17685_3840.n62 103.649
R612 a_17685_3840.n63 a_17685_3840.n31 83.404
R613 a_17685_3840.n31 a_17685_3840.t5 81.437
R614 a_17685_3840.n30 a_17685_3840.n29 73.313
R615 a_17685_3840.n30 a_17685_3840.t4 69.863
R616 a_17685_3840.n29 a_17685_3840.t10 69.653
R617 a_17685_3840.n0 a_17685_3840.n63 66.545
R618 a_17685_3840.n62 a_17685_3840.n61 47.861
R619 a_17685_3840.n24 a_17685_3840.n23 45.936
R620 a_17685_3840.n28 a_17685_3840.n24 41.108
R621 a_17685_3840.n61 a_17685_3840.n55 41.07
R622 a_17685_3840.n31 a_17685_3840.n30 40.307
R623 a_17685_3840.n0 a_17685_3840.t3 29.277
R624 a_17685_3840.t1 a_17685_3840.n0 28.576
R625 a_17685_3840.n0 a_17685_3840.t2 28.565
R626 a_17685_3840.n54 a_17685_3840.n42 24.999
R627 a_17685_3840.n23 a_17685_3840.n11 24.399
R628 a_17685_3840.n32 a_17685_3840.t46 23.529
R629 a_17685_3840.n1 a_17685_3840.t39 23.485
R630 a_17685_3840.n12 a_17685_3840.t31 23.474
R631 a_17685_3840.n43 a_17685_3840.t55 23.456
R632 a_17685_3840.n42 a_17685_3840.t35 15.401
R633 a_17685_3840.n11 a_17685_3840.t50 15.374
R634 a_17685_3840.n53 a_17685_3840.t22 15.341
R635 a_17685_3840.n22 a_17685_3840.t23 15.334
R636 a_17685_3840.n23 a_17685_3840.n22 12.228
R637 a_17685_3840.n54 a_17685_3840.n53 11.433
R638 a_17685_3840.n41 a_17685_3840.n40 10.674
R639 a_17685_3840.n40 a_17685_3840.n39 10.674
R640 a_17685_3840.n39 a_17685_3840.n38 10.674
R641 a_17685_3840.n38 a_17685_3840.n37 10.674
R642 a_17685_3840.n37 a_17685_3840.n36 10.674
R643 a_17685_3840.n36 a_17685_3840.n35 10.674
R644 a_17685_3840.n35 a_17685_3840.n34 10.674
R645 a_17685_3840.n34 a_17685_3840.n33 10.674
R646 a_17685_3840.n33 a_17685_3840.n32 10.674
R647 a_17685_3840.n21 a_17685_3840.n20 10.655
R648 a_17685_3840.n20 a_17685_3840.n19 10.655
R649 a_17685_3840.n19 a_17685_3840.n18 10.655
R650 a_17685_3840.n18 a_17685_3840.n17 10.655
R651 a_17685_3840.n17 a_17685_3840.n16 10.655
R652 a_17685_3840.n16 a_17685_3840.n15 10.655
R653 a_17685_3840.n15 a_17685_3840.n14 10.655
R654 a_17685_3840.n14 a_17685_3840.n13 10.655
R655 a_17685_3840.n13 a_17685_3840.n12 10.655
R656 a_17685_3840.n10 a_17685_3840.n9 10.637
R657 a_17685_3840.n9 a_17685_3840.n8 10.637
R658 a_17685_3840.n8 a_17685_3840.n7 10.637
R659 a_17685_3840.n7 a_17685_3840.n6 10.637
R660 a_17685_3840.n6 a_17685_3840.n5 10.637
R661 a_17685_3840.n5 a_17685_3840.n4 10.637
R662 a_17685_3840.n4 a_17685_3840.n3 10.637
R663 a_17685_3840.n3 a_17685_3840.n2 10.637
R664 a_17685_3840.n2 a_17685_3840.n1 10.637
R665 a_17685_3840.n52 a_17685_3840.n51 10.625
R666 a_17685_3840.n51 a_17685_3840.n50 10.625
R667 a_17685_3840.n50 a_17685_3840.n49 10.625
R668 a_17685_3840.n49 a_17685_3840.n48 10.625
R669 a_17685_3840.n48 a_17685_3840.n47 10.625
R670 a_17685_3840.n47 a_17685_3840.n46 10.625
R671 a_17685_3840.n46 a_17685_3840.n45 10.625
R672 a_17685_3840.n45 a_17685_3840.n44 10.625
R673 a_17685_3840.n44 a_17685_3840.n43 10.625
R674 a_17685_3840.n43 a_17685_3840.t15 8.716
R675 a_17685_3840.n44 a_17685_3840.t21 8.716
R676 a_17685_3840.n45 a_17685_3840.t30 8.716
R677 a_17685_3840.n46 a_17685_3840.t36 8.716
R678 a_17685_3840.n47 a_17685_3840.t13 8.716
R679 a_17685_3840.n48 a_17685_3840.t19 8.716
R680 a_17685_3840.n49 a_17685_3840.t28 8.716
R681 a_17685_3840.n50 a_17685_3840.t26 8.716
R682 a_17685_3840.n51 a_17685_3840.t33 8.716
R683 a_17685_3840.n52 a_17685_3840.t41 8.716
R684 a_17685_3840.n1 a_17685_3840.t47 8.713
R685 a_17685_3840.n2 a_17685_3840.t52 8.713
R686 a_17685_3840.n3 a_17685_3840.t60 8.713
R687 a_17685_3840.n4 a_17685_3840.t16 8.713
R688 a_17685_3840.n5 a_17685_3840.t44 8.713
R689 a_17685_3840.n6 a_17685_3840.t49 8.713
R690 a_17685_3840.n7 a_17685_3840.t56 8.713
R691 a_17685_3840.n8 a_17685_3840.t54 8.713
R692 a_17685_3840.n9 a_17685_3840.t59 8.713
R693 a_17685_3840.n10 a_17685_3840.t18 8.713
R694 a_17685_3840.n12 a_17685_3840.t38 8.708
R695 a_17685_3840.n13 a_17685_3840.t45 8.708
R696 a_17685_3840.n14 a_17685_3840.t51 8.708
R697 a_17685_3840.n15 a_17685_3840.t57 8.708
R698 a_17685_3840.n16 a_17685_3840.t14 8.708
R699 a_17685_3840.n17 a_17685_3840.t20 8.708
R700 a_17685_3840.n18 a_17685_3840.t29 8.708
R701 a_17685_3840.n19 a_17685_3840.t27 8.708
R702 a_17685_3840.n20 a_17685_3840.t34 8.708
R703 a_17685_3840.n21 a_17685_3840.t42 8.708
R704 a_17685_3840.n41 a_17685_3840.t48 8.704
R705 a_17685_3840.n32 a_17685_3840.t53 8.704
R706 a_17685_3840.n33 a_17685_3840.t58 8.704
R707 a_17685_3840.n34 a_17685_3840.t17 8.704
R708 a_17685_3840.n35 a_17685_3840.t24 8.704
R709 a_17685_3840.n36 a_17685_3840.t25 8.704
R710 a_17685_3840.n37 a_17685_3840.t32 8.704
R711 a_17685_3840.n38 a_17685_3840.t40 8.704
R712 a_17685_3840.n39 a_17685_3840.t37 8.704
R713 a_17685_3840.n40 a_17685_3840.t43 8.704
R714 a_17685_3840.n22 a_17685_3840.n21 8.14
R715 a_17685_3840.n42 a_17685_3840.n41 8.128
R716 a_17685_3840.n53 a_17685_3840.n52 8.116
R717 a_17685_3840.n11 a_17685_3840.n10 8.112
R718 a_14266_8900.t16 a_14266_8900.t25 1273.78
R719 a_14266_8900.n3 a_14266_8900.t54 193.916
R720 a_14266_8900.t54 a_14266_8900.t21 113.753
R721 a_14266_8900.t54 a_14266_8900.t11 113.753
R722 a_14266_8900.t54 a_14266_8900.t32 113.753
R723 a_14266_8900.t54 a_14266_8900.t41 113.753
R724 a_14266_8900.t54 a_14266_8900.t52 113.753
R725 a_14266_8900.t54 a_14266_8900.t50 113.753
R726 a_14266_8900.t54 a_14266_8900.t59 113.753
R727 a_14266_8900.t54 a_14266_8900.t18 113.753
R728 a_14266_8900.n2 a_14266_8900.t8 113.753
R729 a_14266_8900.n2 a_14266_8900.t48 113.753
R730 a_14266_8900.n2 a_14266_8900.t42 113.753
R731 a_14266_8900.n2 a_14266_8900.t55 113.753
R732 a_14266_8900.n0 a_14266_8900.t17 113.753
R733 a_14266_8900.n0 a_14266_8900.t34 113.753
R734 a_14266_8900.n1 a_14266_8900.t45 113.753
R735 a_14266_8900.n1 a_14266_8900.t39 113.753
R736 a_14266_8900.n1 a_14266_8900.t13 113.753
R737 a_14266_8900.n1 a_14266_8900.t5 113.753
R738 a_14266_8900.n1 a_14266_8900.t29 113.753
R739 a_14266_8900.n0 a_14266_8900.t23 113.753
R740 a_14266_8900.n0 a_14266_8900.t53 113.753
R741 a_14266_8900.n0 a_14266_8900.t51 113.753
R742 a_14266_8900.n0 a_14266_8900.t60 113.753
R743 a_14266_8900.t47 a_14266_8900.t20 113.753
R744 a_14266_8900.t47 a_14266_8900.t9 113.753
R745 a_14266_8900.t47 a_14266_8900.t49 113.753
R746 a_14266_8900.t47 a_14266_8900.t43 113.753
R747 a_14266_8900.t47 a_14266_8900.t56 113.753
R748 a_14266_8900.n0 a_14266_8900.t19 113.753
R749 a_14266_8900.t47 a_14266_8900.t35 113.753
R750 a_14266_8900.t47 a_14266_8900.t46 113.753
R751 a_14266_8900.t47 a_14266_8900.t40 113.753
R752 a_14266_8900.t47 a_14266_8900.t14 113.753
R753 a_14266_8900.t47 a_14266_8900.t6 113.753
R754 a_14266_8900.t47 a_14266_8900.t30 113.753
R755 a_14266_8900.n0 a_14266_8900.t24 113.753
R756 a_14266_8900.n0 a_14266_8900.t2 113.753
R757 a_14266_8900.n0 a_14266_8900.t61 113.753
R758 a_14266_8900.t47 a_14266_8900.t27 113.753
R759 a_14266_8900.t47 a_14266_8900.t36 113.753
R760 a_14266_8900.t47 a_14266_8900.t31 113.753
R761 a_14266_8900.t47 a_14266_8900.t58 113.753
R762 a_14266_8900.t47 a_14266_8900.t57 113.753
R763 a_14266_8900.t47 a_14266_8900.t7 113.753
R764 a_14266_8900.t54 a_14266_8900.t22 113.753
R765 a_14266_8900.t54 a_14266_8900.t15 113.753
R766 a_14266_8900.t54 a_14266_8900.t33 113.753
R767 a_14266_8900.t54 a_14266_8900.t44 113.753
R768 a_14266_8900.t47 a_14266_8900.t38 113.753
R769 a_14266_8900.t47 a_14266_8900.t12 113.753
R770 a_14266_8900.t47 a_14266_8900.t4 113.753
R771 a_14266_8900.t47 a_14266_8900.t28 113.753
R772 a_14266_8900.t54 a_14266_8900.t37 113.753
R773 a_14266_8900.t54 a_14266_8900.t10 113.753
R774 a_14266_8900.t54 a_14266_8900.t3 113.753
R775 a_14266_8900.t54 a_14266_8900.t26 113.753
R776 a_14266_8900.t1 a_14266_8900.n4 57.619
R777 a_14266_8900.n4 a_14266_8900.n3 43.122
R778 a_14266_8900.n3 a_14266_8900.t0 28.571
R779 a_14266_8900.n4 a_14266_8900.t16 10.022
R780 a_14266_8900.t54 a_14266_8900.n0 5.834
R781 a_14266_8900.t47 a_14266_8900.n1 2.869
R782 a_14266_8900.t54 a_14266_8900.t47 2.813
R783 a_14266_8900.t47 a_14266_8900.n2 2.586
R784 vbiasob.n2 vbiasob.t0 68.426
R785 vbiasob.n0 vbiasob.t3 61.399
R786 vbiasob.n0 vbiasob.t4 60.299
R787 vbiasob.n1 vbiasob.t2 18.573
R788 vbiasob.n3 vbiasob.n2 15.528
R789 vbiasob.n1 vbiasob.t1 5.717
R790 vbiasob.n2 vbiasob.n1 1.006
R791 vbiasob.n3 vbiasob.n0 0.614
R792 vbiasob vbiasob.n3 0.484
R793 a_54432_7362.t0 a_54432_7362.t1 184.898
R794 a_52052_20860.t18 a_52052_20860.n16 2527.24
R795 a_52052_20860.n8 a_52052_20860.t7 212.622
R796 a_52052_20860.n5 a_52052_20860.t16 212.622
R797 a_52052_20860.n12 a_52052_20860.n10 208.271
R798 a_52052_20860.n2 a_52052_20860.n0 208.271
R799 a_52052_20860.n14 a_52052_20860.n12 208.271
R800 a_52052_20860.n9 a_52052_20860.n8 208.271
R801 a_52052_20860.n4 a_52052_20860.n2 208.271
R802 a_52052_20860.n6 a_52052_20860.n5 208.271
R803 a_52052_20860.n7 a_52052_20860.n6 122.265
R804 a_52052_20860.n15 a_52052_20860.n14 121.297
R805 a_52052_20860.n7 a_52052_20860.n4 63.478
R806 a_52052_20860.n15 a_52052_20860.n9 63.217
R807 a_52052_20860.n16 a_52052_20860.n7 38.746
R808 a_52052_20860.n16 a_52052_20860.n15 15.694
R809 a_52052_20860.n8 a_52052_20860.t4 4.351
R810 a_52052_20860.n9 a_52052_20860.t1 4.351
R811 a_52052_20860.n5 a_52052_20860.t13 4.351
R812 a_52052_20860.n6 a_52052_20860.t10 4.351
R813 a_52052_20860.n10 a_52052_20860.t3 4.35
R814 a_52052_20860.n10 a_52052_20860.t8 4.35
R815 a_52052_20860.n11 a_52052_20860.t0 4.35
R816 a_52052_20860.n11 a_52052_20860.t6 4.35
R817 a_52052_20860.n13 a_52052_20860.t5 4.35
R818 a_52052_20860.n13 a_52052_20860.t2 4.35
R819 a_52052_20860.n0 a_52052_20860.t12 4.35
R820 a_52052_20860.n0 a_52052_20860.t17 4.35
R821 a_52052_20860.n1 a_52052_20860.t9 4.35
R822 a_52052_20860.n1 a_52052_20860.t15 4.35
R823 a_52052_20860.n3 a_52052_20860.t14 4.35
R824 a_52052_20860.n3 a_52052_20860.t11 4.35
R825 a_52052_20860.n14 a_52052_20860.n13 0.001
R826 a_52052_20860.n12 a_52052_20860.n11 0.001
R827 a_52052_20860.n4 a_52052_20860.n3 0.001
R828 a_52052_20860.n2 a_52052_20860.n1 0.001
R829 a_56334_20860.n0 a_56334_20860.t1 171.564
R830 a_56334_20860.n0 a_56334_20860.t2 171.563
R831 a_56334_20860.t0 a_56334_20860.n0 171.52
R832 a_23156_5032.n0 a_23156_5032.t7 365.308
R833 a_23156_5032.n4 a_23156_5032.t2 93.107
R834 a_23156_5032.n5 a_23156_5032.n4 75.71
R835 a_23156_5032.n3 a_23156_5032.n2 75.707
R836 a_23156_5032.n2 a_23156_5032.n1 75.707
R837 a_23156_5032.n1 a_23156_5032.n0 75.707
R838 a_23156_5032.n5 a_23156_5032.n3 75.706
R839 a_23156_5032.t6 a_23156_5032.n5 17.401
R840 a_23156_5032.n0 a_23156_5032.t3 17.401
R841 a_23156_5032.n1 a_23156_5032.t0 17.401
R842 a_23156_5032.n2 a_23156_5032.t5 17.401
R843 a_23156_5032.n3 a_23156_5032.t1 17.401
R844 a_23156_5032.n4 a_23156_5032.t4 17.401
R845 a_23436_16644.t46 a_23436_16644.t43 1273.78
R846 a_23436_16644.n3 a_23436_16644.t1 1158.7
R847 a_23436_16644.n3 a_23436_16644.t60 169.095
R848 a_23436_16644.t60 a_23436_16644.t45 113.753
R849 a_23436_16644.t60 a_23436_16644.t5 113.753
R850 a_23436_16644.t60 a_23436_16644.t21 113.753
R851 a_23436_16644.t60 a_23436_16644.t20 113.753
R852 a_23436_16644.t60 a_23436_16644.t2 113.753
R853 a_23436_16644.t60 a_23436_16644.t17 113.753
R854 a_23436_16644.t60 a_23436_16644.t37 113.753
R855 a_23436_16644.t60 a_23436_16644.t33 113.753
R856 a_23436_16644.n2 a_23436_16644.t44 113.753
R857 a_23436_16644.n2 a_23436_16644.t59 113.753
R858 a_23436_16644.n2 a_23436_16644.t14 113.753
R859 a_23436_16644.n2 a_23436_16644.t32 113.753
R860 a_23436_16644.n0 a_23436_16644.t10 113.753
R861 a_23436_16644.n0 a_23436_16644.t28 113.753
R862 a_23436_16644.n1 a_23436_16644.t26 113.753
R863 a_23436_16644.n1 a_23436_16644.t34 113.753
R864 a_23436_16644.n1 a_23436_16644.t47 113.753
R865 a_23436_16644.n1 a_23436_16644.t6 113.753
R866 a_23436_16644.n1 a_23436_16644.t24 113.753
R867 a_23436_16644.n0 a_23436_16644.t50 113.753
R868 a_23436_16644.n0 a_23436_16644.t22 113.753
R869 a_23436_16644.n0 a_23436_16644.t40 113.753
R870 a_23436_16644.n0 a_23436_16644.t58 113.753
R871 a_23436_16644.t12 a_23436_16644.t56 113.753
R872 a_23436_16644.t12 a_23436_16644.t8 113.753
R873 a_23436_16644.t12 a_23436_16644.t18 113.753
R874 a_23436_16644.t12 a_23436_16644.t38 113.753
R875 a_23436_16644.t12 a_23436_16644.t54 113.753
R876 a_23436_16644.n0 a_23436_16644.t11 113.753
R877 a_23436_16644.t12 a_23436_16644.t29 113.753
R878 a_23436_16644.t12 a_23436_16644.t27 113.753
R879 a_23436_16644.t12 a_23436_16644.t35 113.753
R880 a_23436_16644.t12 a_23436_16644.t48 113.753
R881 a_23436_16644.t12 a_23436_16644.t7 113.753
R882 a_23436_16644.t12 a_23436_16644.t25 113.753
R883 a_23436_16644.n0 a_23436_16644.t51 113.753
R884 a_23436_16644.n0 a_23436_16644.t23 113.753
R885 a_23436_16644.n0 a_23436_16644.t41 113.753
R886 a_23436_16644.t12 a_23436_16644.t61 113.753
R887 a_23436_16644.t12 a_23436_16644.t57 113.753
R888 a_23436_16644.t12 a_23436_16644.t9 113.753
R889 a_23436_16644.t12 a_23436_16644.t19 113.753
R890 a_23436_16644.t12 a_23436_16644.t39 113.753
R891 a_23436_16644.t12 a_23436_16644.t55 113.753
R892 a_23436_16644.t60 a_23436_16644.t15 113.753
R893 a_23436_16644.t60 a_23436_16644.t36 113.753
R894 a_23436_16644.t60 a_23436_16644.t53 113.753
R895 a_23436_16644.t60 a_23436_16644.t52 113.753
R896 a_23436_16644.t12 a_23436_16644.t4 113.753
R897 a_23436_16644.t12 a_23436_16644.t13 113.753
R898 a_23436_16644.t12 a_23436_16644.t31 113.753
R899 a_23436_16644.t12 a_23436_16644.t49 113.753
R900 a_23436_16644.t60 a_23436_16644.t30 113.753
R901 a_23436_16644.t60 a_23436_16644.t42 113.753
R902 a_23436_16644.t60 a_23436_16644.t3 113.753
R903 a_23436_16644.t60 a_23436_16644.t16 113.753
R904 a_23436_16644.t0 a_23436_16644.n3 59.624
R905 a_23436_16644.t60 a_23436_16644.t46 6.578
R906 a_23436_16644.t60 a_23436_16644.n0 5.834
R907 a_23436_16644.t12 a_23436_16644.n1 2.869
R908 a_23436_16644.t12 a_23436_16644.n2 2.586
R909 a_23436_16644.t60 a_23436_16644.t12 2.576
R910 a_25778_4988.n0 a_25778_4988.t7 334.707
R911 a_25778_4988.n4 a_25778_4988.t2 93.107
R912 a_25778_4988.n5 a_25778_4988.n4 75.71
R913 a_25778_4988.n3 a_25778_4988.n2 75.707
R914 a_25778_4988.n2 a_25778_4988.n1 75.707
R915 a_25778_4988.n1 a_25778_4988.n0 75.707
R916 a_25778_4988.n5 a_25778_4988.n3 75.706
R917 a_25778_4988.t6 a_25778_4988.n5 17.401
R918 a_25778_4988.n0 a_25778_4988.t3 17.401
R919 a_25778_4988.n1 a_25778_4988.t0 17.401
R920 a_25778_4988.n2 a_25778_4988.t5 17.401
R921 a_25778_4988.n3 a_25778_4988.t1 17.401
R922 a_25778_4988.n4 a_25778_4988.t4 17.401
R923 a_22429_17162.t34 a_22429_17162.t11 1273.78
R924 a_22429_17162.n3 a_22429_17162.t34 132.569
R925 a_22429_17162.t29 a_22429_17162.t13 113.753
R926 a_22429_17162.t29 a_22429_17162.t7 113.753
R927 a_22429_17162.t29 a_22429_17162.t31 113.753
R928 a_22429_17162.t29 a_22429_17162.t39 113.753
R929 a_22429_17162.t29 a_22429_17162.t30 113.753
R930 a_22429_17162.t29 a_22429_17162.t28 113.753
R931 a_22429_17162.t29 a_22429_17162.t44 113.753
R932 a_22429_17162.t29 a_22429_17162.t58 113.753
R933 a_22429_17162.n2 a_22429_17162.t57 113.753
R934 a_22429_17162.n2 a_22429_17162.t27 113.753
R935 a_22429_17162.n2 a_22429_17162.t24 113.753
R936 a_22429_17162.n2 a_22429_17162.t36 113.753
R937 a_22429_17162.n0 a_22429_17162.t17 113.753
R938 a_22429_17162.n0 a_22429_17162.t33 113.753
R939 a_22429_17162.n1 a_22429_17162.t47 113.753
R940 a_22429_17162.n1 a_22429_17162.t40 113.753
R941 a_22429_17162.n1 a_22429_17162.t15 113.753
R942 a_22429_17162.n1 a_22429_17162.t9 113.753
R943 a_22429_17162.n1 a_22429_17162.t25 113.753
R944 a_22429_17162.n0 a_22429_17162.t21 113.753
R945 a_22429_17162.n0 a_22429_17162.t54 113.753
R946 a_22429_17162.n0 a_22429_17162.t52 113.753
R947 a_22429_17162.n0 a_22429_17162.t2 113.753
R948 a_22429_17162.n1 a_22429_17162.t19 113.753
R949 a_22429_17162.n1 a_22429_17162.t12 113.753
R950 a_22429_17162.n1 a_22429_17162.t50 113.753
R951 a_22429_17162.n1 a_22429_17162.t45 113.753
R952 a_22429_17162.n1 a_22429_17162.t59 113.753
R953 a_22429_17162.n0 a_22429_17162.t18 113.753
R954 a_22429_17162.n1 a_22429_17162.t35 113.753
R955 a_22429_17162.n1 a_22429_17162.t48 113.753
R956 a_22429_17162.n1 a_22429_17162.t41 113.753
R957 a_22429_17162.n1 a_22429_17162.t16 113.753
R958 a_22429_17162.n1 a_22429_17162.t10 113.753
R959 a_22429_17162.n1 a_22429_17162.t26 113.753
R960 a_22429_17162.n0 a_22429_17162.t22 113.753
R961 a_22429_17162.n0 a_22429_17162.t55 113.753
R962 a_22429_17162.n0 a_22429_17162.t53 113.753
R963 a_22429_17162.n1 a_22429_17162.t3 113.753
R964 a_22429_17162.n1 a_22429_17162.t20 113.753
R965 a_22429_17162.n1 a_22429_17162.t14 113.753
R966 a_22429_17162.n1 a_22429_17162.t51 113.753
R967 a_22429_17162.n1 a_22429_17162.t46 113.753
R968 a_22429_17162.n1 a_22429_17162.t60 113.753
R969 a_22429_17162.t29 a_22429_17162.t49 113.753
R970 a_22429_17162.t29 a_22429_17162.t43 113.753
R971 a_22429_17162.t29 a_22429_17162.t61 113.753
R972 a_22429_17162.t29 a_22429_17162.t8 113.753
R973 a_22429_17162.n1 a_22429_17162.t5 113.753
R974 a_22429_17162.n1 a_22429_17162.t42 113.753
R975 a_22429_17162.n1 a_22429_17162.t38 113.753
R976 a_22429_17162.n1 a_22429_17162.t56 113.753
R977 a_22429_17162.t29 a_22429_17162.t37 113.753
R978 a_22429_17162.t29 a_22429_17162.t6 113.753
R979 a_22429_17162.t29 a_22429_17162.t4 113.753
R980 a_22429_17162.t29 a_22429_17162.t23 113.753
R981 a_22429_17162.t1 a_22429_17162.n3 77.367
R982 a_22429_17162.n3 a_22429_17162.t0 28.578
R983 a_22429_17162.t29 a_22429_17162.n0 5.834
R984 a_22429_17162.t34 a_22429_17162.t29 5.391
R985 a_22429_17162.n1 a_22429_17162.n2 4.056
R986 a_22429_17162.n1 a_22429_17162.t32 2.864
R987 a_22429_17162.t29 a_22429_17162.n1 2.813
R988 a_56272_15934.t1 a_56272_15934.t0 409.924
R989 a_49858_3690.n0 a_49858_3690.t7 19.742
R990 a_49858_3690.n0 a_49858_3690.t5 18.733
R991 a_49858_3690.t2 a_49858_3690.n1 18.498
R992 a_49858_3690.n3 a_49858_3690.t3 17.928
R993 a_49858_3690.n0 a_49858_3690.t8 16.208
R994 a_49858_3690.n1 a_49858_3690.t1 15.946
R995 a_49858_3690.n2 a_49858_3690.t10 9.868
R996 a_49858_3690.n2 a_49858_3690.t6 7.325
R997 a_49858_3690.n2 a_49858_3690.t11 6.179
R998 a_49858_3690.n1 a_49858_3690.t0 5.514
R999 a_49858_3690.n0 a_49858_3690.t12 5.514
R1000 a_49858_3690.n3 a_49858_3690.t4 5.512
R1001 a_49858_3690.n1 a_49858_3690.n0 4.479
R1002 a_49858_3690.n4 a_49858_3690.n3 4.094
R1003 a_49858_3690.n4 a_49858_3690.t9 3.856
R1004 a_49858_3690.n0 a_49858_3690.n4 3.301
R1005 a_49858_3690.n0 a_49858_3690.n2 2.265
R1006 a_49916_3664.t1 a_49916_3664.t2 33.597
R1007 a_49916_3664.t0 a_49916_3664.t1 13.614
R1008 a_49916_3664.t1 a_49916_3664.t3 11.692
R1009 a_28578_5014.n5 a_28578_5014.t7 265.844
R1010 a_28578_5014.n0 a_28578_5014.t5 93.107
R1011 a_28578_5014.n5 a_28578_5014.n4 75.71
R1012 a_28578_5014.n1 a_28578_5014.n0 75.707
R1013 a_28578_5014.n2 a_28578_5014.n1 75.707
R1014 a_28578_5014.n3 a_28578_5014.n2 75.707
R1015 a_28578_5014.n4 a_28578_5014.n3 75.707
R1016 a_28578_5014.t6 a_28578_5014.n5 17.401
R1017 a_28578_5014.n4 a_28578_5014.t3 17.401
R1018 a_28578_5014.n3 a_28578_5014.t1 17.401
R1019 a_28578_5014.n2 a_28578_5014.t4 17.401
R1020 a_28578_5014.n1 a_28578_5014.t2 17.401
R1021 a_28578_5014.n0 a_28578_5014.t0 17.401
R1022 a_51516_3690.n1 a_51516_3690.t3 19.231
R1023 a_51516_3690.n0 a_51516_3690.t2 17.234
R1024 a_51516_3690.n2 a_51516_3690.t4 14.994
R1025 a_51516_3690.n0 a_51516_3690.t1 14.151
R1026 a_51516_3690.n1 a_51516_3690.t5 13.856
R1027 a_51516_3690.t0 a_51516_3690.n0 7.827
R1028 a_51516_3690.n1 a_51516_3690.n2 5.632
R1029 a_51516_3690.n2 a_51516_3690.t6 3.653
R1030 a_51516_3690.n0 a_51516_3690.n1 3.447
R1031 a_50583_13108.n0 a_50583_13108.t1 1776.66
R1032 a_50583_13108.n0 a_50583_13108.t2 171.607
R1033 a_50583_13108.t0 a_50583_13108.n0 171.607
R1034 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n4 1158.04
R1035 Fvco_By4_QPH_bar.t10 Fvco_By4_QPH_bar.t9 731.89
R1036 Fvco_By4_QPH_bar.t5 Fvco_By4_QPH_bar.t14 719.978
R1037 Fvco_By4_QPH_bar.t8 Fvco_By4_QPH_bar.t18 710.965
R1038 Fvco_By4_QPH_bar.t7 Fvco_By4_QPH_bar.t19 710.965
R1039 Fvco_By4_QPH_bar.t6 Fvco_By4_QPH_bar.t13 710.965
R1040 Fvco_By4_QPH_bar.t18 Fvco_By4_QPH_bar.t17 579.889
R1041 Fvco_By4_QPH_bar.t19 Fvco_By4_QPH_bar.t15 579.889
R1042 Fvco_By4_QPH_bar.t13 Fvco_By4_QPH_bar.t12 579.889
R1043 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.t7 570.03
R1044 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.t6 563.963
R1045 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.t8 557.83
R1046 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n2 458.46
R1047 Fvco_By4_QPH_bar.n8 Fvco_By4_QPH_bar.n7 435.858
R1048 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.t16 417.917
R1049 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.t11 414.213
R1050 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.t4 414.167
R1051 Fvco_By4_QPH_bar.n8 Fvco_By4_QPH_bar.t5 245.573
R1052 Fvco_By4_QPH_bar.n9 Fvco_By4_QPH_bar.t10 244.389
R1053 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n9 188.615
R1054 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.n6 149.023
R1055 Fvco_By4_QPH_bar.n9 Fvco_By4_QPH_bar.n8 130.017
R1056 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.n3 50.411
R1057 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.n1 24.956
R1058 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.n0 24.185
R1059 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t1 21.888
R1060 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t0 21.888
R1061 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t2 20
R1062 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t3 20
R1063 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.n5 1.452
R1064 a_27762_11446.t11 a_27762_11446.t48 1273.78
R1065 a_27762_11446.t47 a_27762_11446.t13 113.753
R1066 a_27762_11446.t47 a_27762_11446.t23 113.753
R1067 a_27762_11446.t47 a_27762_11446.t39 113.753
R1068 a_27762_11446.t47 a_27762_11446.t56 113.753
R1069 a_27762_11446.t47 a_27762_11446.t45 113.753
R1070 a_27762_11446.t47 a_27762_11446.t60 113.753
R1071 a_27762_11446.t47 a_27762_11446.t9 113.753
R1072 a_27762_11446.t47 a_27762_11446.t30 113.753
R1073 a_27762_11446.n2 a_27762_11446.t25 113.753
R1074 a_27762_11446.n2 a_27762_11446.t37 113.753
R1075 a_27762_11446.n2 a_27762_11446.t53 113.753
R1076 a_27762_11446.n2 a_27762_11446.t7 113.753
R1077 a_27762_11446.n0 a_27762_11446.t28 113.753
R1078 a_27762_11446.n0 a_27762_11446.t41 113.753
R1079 a_27762_11446.n1 a_27762_11446.t58 113.753
R1080 a_27762_11446.n1 a_27762_11446.t51 113.753
R1081 a_27762_11446.n1 a_27762_11446.t5 113.753
R1082 a_27762_11446.n1 a_27762_11446.t20 113.753
R1083 a_27762_11446.n1 a_27762_11446.t35 113.753
R1084 a_27762_11446.n0 a_27762_11446.t15 113.753
R1085 a_27762_11446.n0 a_27762_11446.t46 113.753
R1086 a_27762_11446.n0 a_27762_11446.t61 113.753
R1087 a_27762_11446.n0 a_27762_11446.t10 113.753
R1088 a_27762_11446.t21 a_27762_11446.t31 113.753
R1089 a_27762_11446.t21 a_27762_11446.t26 113.753
R1090 a_27762_11446.t21 a_27762_11446.t38 113.753
R1091 a_27762_11446.t21 a_27762_11446.t54 113.753
R1092 a_27762_11446.t21 a_27762_11446.t8 113.753
R1093 a_27762_11446.n0 a_27762_11446.t29 113.753
R1094 a_27762_11446.t21 a_27762_11446.t42 113.753
R1095 a_27762_11446.t21 a_27762_11446.t59 113.753
R1096 a_27762_11446.t21 a_27762_11446.t52 113.753
R1097 a_27762_11446.t21 a_27762_11446.t6 113.753
R1098 a_27762_11446.t21 a_27762_11446.t22 113.753
R1099 a_27762_11446.t21 a_27762_11446.t36 113.753
R1100 a_27762_11446.n0 a_27762_11446.t16 113.753
R1101 a_27762_11446.n0 a_27762_11446.t3 113.753
R1102 a_27762_11446.n0 a_27762_11446.t17 113.753
R1103 a_27762_11446.t21 a_27762_11446.t32 113.753
R1104 a_27762_11446.t21 a_27762_11446.t44 113.753
R1105 a_27762_11446.t21 a_27762_11446.t43 113.753
R1106 a_27762_11446.t21 a_27762_11446.t55 113.753
R1107 a_27762_11446.t21 a_27762_11446.t12 113.753
R1108 a_27762_11446.t21 a_27762_11446.t24 113.753
R1109 a_27762_11446.t47 a_27762_11446.t14 113.753
R1110 a_27762_11446.t47 a_27762_11446.t27 113.753
R1111 a_27762_11446.t47 a_27762_11446.t40 113.753
R1112 a_27762_11446.t47 a_27762_11446.t57 113.753
R1113 a_27762_11446.t21 a_27762_11446.t50 113.753
R1114 a_27762_11446.t21 a_27762_11446.t4 113.753
R1115 a_27762_11446.t21 a_27762_11446.t19 113.753
R1116 a_27762_11446.t21 a_27762_11446.t34 113.753
R1117 a_27762_11446.t47 a_27762_11446.t49 113.753
R1118 a_27762_11446.t47 a_27762_11446.t2 113.753
R1119 a_27762_11446.t47 a_27762_11446.t18 113.753
R1120 a_27762_11446.t47 a_27762_11446.t33 113.753
R1121 a_27762_11446.n4 a_27762_11446.n3 88.886
R1122 a_27762_11446.n4 a_27762_11446.t0 81.996
R1123 a_27762_11446.t1 a_27762_11446.n4 59.267
R1124 a_27762_11446.t47 a_27762_11446.n0 5.834
R1125 a_27762_11446.n3 a_27762_11446.t11 4.994
R1126 a_27762_11446.n3 a_27762_11446.t47 4.809
R1127 a_27762_11446.t21 a_27762_11446.n1 2.869
R1128 a_27762_11446.t47 a_27762_11446.t21 2.8
R1129 a_27762_11446.t21 a_27762_11446.n2 2.586
R1130 a_44752_16348.t2 a_44752_16348.n2 349.137
R1131 a_44752_16348.n1 a_44752_16348.t1 197.553
R1132 a_44752_16348.n0 a_44752_16348.t3 178.539
R1133 a_44752_16348.n0 a_44752_16348.t4 122.603
R1134 a_44752_16348.n1 a_44752_16348.t0 114.713
R1135 a_44752_16348.n2 a_44752_16348.n0 95.215
R1136 a_44752_16348.n2 a_44752_16348.n1 26.034
R1137 a_51138_19904.t0 a_51138_19904.n0 171.568
R1138 a_51138_19904.n0 a_51138_19904.t1 171.564
R1139 a_51138_19904.n0 a_51138_19904.t2 171.52
R1140 a_14832_12082.n1 a_14832_12082.t3 434.515
R1141 a_14832_12082.n0 a_14832_12082.t2 217.163
R1142 a_14832_12082.t0 a_14832_12082.n1 52.152
R1143 a_14832_12082.n0 a_14832_12082.t1 3.106
R1144 a_14832_12082.n1 a_14832_12082.n0 0.908
R1145 a_23160_10936.n0 a_23160_10936.t0 391.966
R1146 a_23160_10936.t6 a_23160_10936.n5 93.107
R1147 a_23160_10936.n1 a_23160_10936.n0 75.707
R1148 a_23160_10936.n5 a_23160_10936.n4 75.707
R1149 a_23160_10936.n4 a_23160_10936.n3 75.707
R1150 a_23160_10936.n3 a_23160_10936.n2 75.707
R1151 a_23160_10936.n2 a_23160_10936.n1 75.707
R1152 a_23160_10936.n0 a_23160_10936.t7 17.401
R1153 a_23160_10936.n1 a_23160_10936.t3 17.401
R1154 a_23160_10936.n2 a_23160_10936.t1 17.401
R1155 a_23160_10936.n3 a_23160_10936.t4 17.401
R1156 a_23160_10936.n4 a_23160_10936.t2 17.401
R1157 a_23160_10936.n5 a_23160_10936.t5 17.401
R1158 a_28438_10874.n0 a_28438_10874.t7 338.927
R1159 a_28438_10874.n4 a_28438_10874.t3 93.107
R1160 a_28438_10874.n5 a_28438_10874.n4 75.71
R1161 a_28438_10874.n1 a_28438_10874.n0 75.708
R1162 a_28438_10874.n3 a_28438_10874.n2 75.707
R1163 a_28438_10874.n2 a_28438_10874.n1 75.707
R1164 a_28438_10874.n5 a_28438_10874.n3 75.706
R1165 a_28438_10874.t6 a_28438_10874.n5 17.401
R1166 a_28438_10874.n0 a_28438_10874.t4 17.401
R1167 a_28438_10874.n1 a_28438_10874.t0 17.401
R1168 a_28438_10874.n2 a_28438_10874.t5 17.401
R1169 a_28438_10874.n3 a_28438_10874.t1 17.401
R1170 a_28438_10874.n4 a_28438_10874.t2 17.401
R1171 a_14910_6932.n1 a_14910_6932.t3 434.494
R1172 a_14910_6932.n0 a_14910_6932.t2 217.163
R1173 a_14910_6932.t0 a_14910_6932.n1 52.318
R1174 a_14910_6932.n0 a_14910_6932.t1 3.106
R1175 a_14910_6932.n1 a_14910_6932.n0 0.906
R1176 a_64603_26128.t6 a_64603_26128.t4 2276.65
R1177 a_64603_26128.n0 a_64603_26128.t5 1000.95
R1178 a_64603_26128.t3 a_64603_26128.n1 779.232
R1179 a_64603_26128.n1 a_64603_26128.t2 589.347
R1180 a_64603_26128.n2 a_64603_26128.t3 560.159
R1181 a_64603_26128.n1 a_64603_26128.n0 298.84
R1182 a_64603_26128.n0 a_64603_26128.t7 176.733
R1183 a_64603_26128.t0 a_64603_26128.n3 135.884
R1184 a_64603_26128.n2 a_64603_26128.t6 124.034
R1185 a_64603_26128.n3 a_64603_26128.t1 62.096
R1186 a_64603_26128.n3 a_64603_26128.n2 33.009
R1187 a_26016_10878.n5 a_26016_10878.t7 305.609
R1188 a_26016_10878.n0 a_26016_10878.t5 93.107
R1189 a_26016_10878.n5 a_26016_10878.n4 75.71
R1190 a_26016_10878.n1 a_26016_10878.n0 75.707
R1191 a_26016_10878.n2 a_26016_10878.n1 75.707
R1192 a_26016_10878.n3 a_26016_10878.n2 75.707
R1193 a_26016_10878.n4 a_26016_10878.n3 75.707
R1194 a_26016_10878.t6 a_26016_10878.n5 17.401
R1195 a_26016_10878.n4 a_26016_10878.t2 17.401
R1196 a_26016_10878.n3 a_26016_10878.t0 17.401
R1197 a_26016_10878.n2 a_26016_10878.t3 17.401
R1198 a_26016_10878.n1 a_26016_10878.t1 17.401
R1199 a_26016_10878.n0 a_26016_10878.t4 17.401
R1200 a_77280_24640.n1 a_77280_24640.t3 263.373
R1201 a_77280_24640.t0 a_77280_24640.n2 61.061
R1202 a_77280_24640.n0 a_77280_24640.t4 14.065
R1203 a_77280_24640.n0 a_77280_24640.t2 4.819
R1204 a_77280_24640.n2 a_77280_24640.n0 2.726
R1205 a_77280_24640.n1 a_77280_24640.t1 1.368
R1206 a_77280_24640.n2 a_77280_24640.n1 0.571
R1207 a_77254_23336.t6 a_77254_23336.n3 95.488
R1208 a_77254_23336.n0 a_77254_23336.t2 52.208
R1209 a_77254_23336.n3 a_77254_23336.n2 13.658
R1210 a_77254_23336.n3 a_77254_23336.t5 4.572
R1211 a_77254_23336.n1 a_77254_23336.t1 3.848
R1212 a_77254_23336.n0 a_77254_23336.t4 1.482
R1213 a_77254_23336.n2 a_77254_23336.n1 1.338
R1214 a_77254_23336.n1 a_77254_23336.t3 0.701
R1215 a_77254_23336.n2 a_77254_23336.n0 0.15
R1216 a_77254_23336.t5 a_77254_23336.t0 0.049
R1217 a_24410_25128.n1 a_24410_25128.t3 434.509
R1218 a_24410_25128.n0 a_24410_25128.t2 217.163
R1219 a_24410_25128.t0 a_24410_25128.n1 52.459
R1220 a_24410_25128.n0 a_24410_25128.t1 3.106
R1221 a_24410_25128.n1 a_24410_25128.n0 0.899
R1222 a_23308_802.n1 a_23308_802.t2 434.515
R1223 a_23308_802.n0 a_23308_802.t3 217.163
R1224 a_23308_802.t0 a_23308_802.n1 52.152
R1225 a_23308_802.n0 a_23308_802.t1 3.106
R1226 a_23308_802.n1 a_23308_802.n0 0.908
R1227 a_57710_5326.n0 a_57710_5326.t1 85.561
R1228 a_57710_5326.n1 a_57710_5326.t3 85.561
R1229 a_57710_5326.n0 a_57710_5326.t5 39.685
R1230 a_57710_5326.n1 a_57710_5326.t0 17.517
R1231 a_57710_5326.t2 a_57710_5326.n3 5.8
R1232 a_57710_5326.n3 a_57710_5326.t4 5.8
R1233 a_57710_5326.n3 a_57710_5326.n2 0.736
R1234 a_57710_5326.n2 a_57710_5326.n0 0.231
R1235 a_57710_5326.n2 a_57710_5326.n1 0.206
R1236 a_32948_24994.n1 a_32948_24994.t3 434.487
R1237 a_32948_24994.n0 a_32948_24994.t2 217.163
R1238 a_32948_24994.t0 a_32948_24994.n1 52.153
R1239 a_32948_24994.n0 a_32948_24994.t1 3.106
R1240 a_32948_24994.n1 a_32948_24994.n0 0.887
R1241 a_28790_25040.n1 a_28790_25040.t3 434.517
R1242 a_28790_25040.n0 a_28790_25040.t2 217.163
R1243 a_28790_25040.t0 a_28790_25040.n1 52.317
R1244 a_28790_25040.n0 a_28790_25040.t1 3.106
R1245 a_28790_25040.n1 a_28790_25040.n0 0.907
R1246 a_50032_16080.t0 a_50032_16080.t1 414.247
R1247 a_50511_16072.n4 a_50511_16072.n3 524.893
R1248 a_50511_16072.n4 a_50511_16072.t8 256.935
R1249 a_50511_16072.t5 a_50511_16072.n1 8.763
R1250 a_50511_16072.n2 a_50511_16072.t0 8.705
R1251 a_50511_16072.n1 a_50511_16072.t1 8.7
R1252 a_50511_16072.n1 a_50511_16072.t2 8.7
R1253 a_50511_16072.n0 a_50511_16072.t3 8.7
R1254 a_50511_16072.n0 a_50511_16072.t4 8.7
R1255 a_50511_16072.n3 a_50511_16072.t7 5.844
R1256 a_50511_16072.n3 a_50511_16072.t6 5.744
R1257 a_50511_16072.t8 a_50511_16072.t9 1.22
R1258 a_50511_16072.n1 a_50511_16072.n0 0.137
R1259 a_50511_16072.n0 a_50511_16072.n2 0.133
R1260 a_50511_16072.n0 a_50511_16072.n4 0.122
R1261 a_38070_8852.n1 a_38070_8852.t3 434.515
R1262 a_38070_8852.n0 a_38070_8852.t2 217.163
R1263 a_38070_8852.t0 a_38070_8852.n1 52.152
R1264 a_38070_8852.n0 a_38070_8852.t1 3.106
R1265 a_38070_8852.n1 a_38070_8852.n0 0.908
R1266 a_30384_802.n1 a_30384_802.t3 434.478
R1267 a_30384_802.n0 a_30384_802.t2 217.163
R1268 a_30384_802.t0 a_30384_802.n1 52.152
R1269 a_30384_802.n0 a_30384_802.t1 3.106
R1270 a_30384_802.n1 a_30384_802.n0 0.885
R1271 a_77598_24640.n1 a_77598_24640.t3 256.234
R1272 a_77598_24640.n0 a_77598_24640.t2 12.058
R1273 a_77598_24640.t0 a_77598_24640.n2 11.463
R1274 a_77598_24640.n0 a_77598_24640.t4 4.624
R1275 a_77598_24640.n1 a_77598_24640.t1 2.155
R1276 a_77598_24640.n2 a_77598_24640.n0 1.194
R1277 a_77598_24640.n2 a_77598_24640.n1 0.952
R1278 a_77572_23336.t4 a_77572_23336.n3 7.523
R1279 a_77572_23336.n0 a_77572_23336.t1 3.01
R1280 a_77572_23336.n1 a_77572_23336.t6 2.635
R1281 a_77572_23336.n2 a_77572_23336.t0 1.86
R1282 a_77572_23336.n3 a_77572_23336.n2 1.672
R1283 a_77572_23336.n3 a_77572_23336.n1 1.093
R1284 a_77572_23336.n0 a_77572_23336.t3 0.778
R1285 a_77572_23336.n2 a_77572_23336.t2 0.727
R1286 a_77572_23336.n1 a_77572_23336.n0 0.166
R1287 a_77572_23336.t6 a_77572_23336.t5 0.037
R1288 a_46856_21176.t0 a_46856_21176.t1 343.213
R1289 a_51138_21494.t1 a_51138_21494.t0 501.405
R1290 vbiasot.t0 vbiasot.t2 17.477
R1291 vbiasot.t0 vbiasot.t1 12.163
R1292 vbiasot vbiasot.t0 10.441
R1293 a_46856_19268.n0 a_46856_19268.t1 2113.41
R1294 a_46856_19268.n0 a_46856_19268.t2 171.607
R1295 a_46856_19268.t0 a_46856_19268.n0 171.607
R1296 vbiasbuffer.n0 vbiasbuffer.t0 137.132
R1297 vbiasbuffer.n2 vbiasbuffer.t4 125.304
R1298 vbiasbuffer.n2 vbiasbuffer.t3 120.586
R1299 vbiasbuffer vbiasbuffer.n1 22.704
R1300 vbiasbuffer.n1 vbiasbuffer.t2 13.427
R1301 vbiasbuffer.n1 vbiasbuffer.n0 8.397
R1302 vbiasbuffer.n0 vbiasbuffer.t1 5.717
R1303 vbiasbuffer vbiasbuffer.n2 0.631
R1304 a_51826_16054.t1 a_51826_16054.t0 445.429
R1305 a_54452_7044.t1 a_54452_7044.t0 178.373
R1306 a_22972_23306.t3 a_22972_23306.n2 172.018
R1307 a_22972_23306.n2 a_22972_23306.t4 171.695
R1308 a_22972_23306.n2 a_22972_23306.n1 73.126
R1309 a_22972_23306.n1 a_22972_23306.t2 28.576
R1310 a_22972_23306.n0 a_22972_23306.t0 28.565
R1311 a_22972_23306.n0 a_22972_23306.t1 28.565
R1312 a_22972_23306.n1 a_22972_23306.n0 3.497
C61 vbiasr gnd 139.20fF $ **FLOATING
C62 vbiasot gnd 36.48fF $ **FLOATING
C63 a_51334_14126# gnd 5.94fF
C64 a_50320_14126# gnd 7.42fF
C65 a_56602_11692# gnd 4.81fF
C66 a_55602_11692# gnd 5.68fF
C67 a_51276_14152# gnd 3.34fF
C68 a_51636_13108# gnd 8.30fF
C69 a_51041_13108# gnd 10.28fF
C70 a_50262_14152# gnd 3.87fF
C71 vbiasob gnd 12.28fF $ **FLOATING
C72 a_47760_15642# gnd 2.83fF
C73 vbiasbuffer gnd 27.30fF $ **FLOATING
C74 a_43010_16058# gnd 4.05fF
C75 a_42782_16060# gnd 4.44fF
C76 a_42574_15624# gnd 5.31fF
C77 a_42550_16062# gnd 4.20fF
C78 a_45810_16322# gnd 24.39fF
C79 a_44810_16322# gnd 24.18fF
C80 Vso8b gnd 20.82fF
C81 Vso7b gnd 14.60fF
C82 a_4226_11420# gnd 8.28fF
C83 a_4288_11534# gnd 5.07fF
C84 a_4226_11612# gnd 7.54fF
C85 a_4288_11726# gnd 6.25fF
C86 a_4226_11804# gnd 7.73fF
C87 Vso5b gnd 7.67fF
C88 Vso4b gnd 47.35fF
C89 Vso6b gnd 5.87fF
C90 a_4288_11918# gnd 5.18fF
C91 a_4226_11996# gnd 8.59fF
C92 a_4288_12110# gnd 6.31fF
C93 v9m gnd 13.79fF
C94 a_4226_12188# gnd 6.34fF
C95 Fvco_By4_QPH_bar gnd 26.88fF $ **FLOATING
C96 Fvco_By4_QPH gnd 36.85fF $ **FLOATING
C97 reset gnd 45.36fF $ **FLOATING
C98 Fvco gnd 124.77fF
C99 Vso3b gnd 26.66fF
C100 Vso2b gnd 21.36fF
C101 Vso1b gnd 22.16fF
C102 vctrl gnd 12.55fF
C103 a_33808_31746# gnd 16.63fF
C104 vinit gnd 191.08fF $ **FLOATING
C105 a_34044_31208# gnd 377.15fF
C106 a_9354_33563# gnd 376.67fF
C107 vdd gnd 6130.32fF
C108 a_22972_23306.n2 gnd 2.07fF $ **FLOATING
C109 a_54452_7044.t0 gnd 2.83fF
C110 vbiasbuffer.n1 gnd 11.83fF $ **FLOATING
C111 a_46856_19268.n0 gnd 7.50fF $ **FLOATING
C112 vbiasot.t0 gnd 8.65fF
C113 a_51138_21494.t0 gnd 2.55fF
C114 a_51138_21494.t1 gnd 3.48fF
C115 a_77572_23336.t1 gnd 72.17fF
C116 a_77572_23336.t3 gnd 49.69fF
C117 a_77572_23336.n0 gnd 52.35fF $ **FLOATING
C118 a_77572_23336.t5 gnd 37.84fF $ **FLOATING
C119 a_77572_23336.t6 gnd 61.50fF $ **FLOATING
C120 a_77572_23336.n1 gnd 84.84fF $ **FLOATING
C121 a_77572_23336.t2 gnd 42.57fF
C122 a_77572_23336.t0 gnd 52.39fF
C123 a_77572_23336.n2 gnd 60.74fF $ **FLOATING
C124 a_77572_23336.n3 gnd 66.26fF $ **FLOATING
C125 a_77598_24640.t2 gnd 44.04fF $ **FLOATING
C126 a_77598_24640.t4 gnd 42.02fF $ **FLOATING
C127 a_77598_24640.n0 gnd 35.23fF $ **FLOATING
C128 a_77598_24640.t3 gnd 70.35fF $ **FLOATING
C129 a_77598_24640.t1 gnd 50.88fF $ **FLOATING
C130 a_77598_24640.n1 gnd 43.65fF $ **FLOATING
C131 a_77598_24640.n2 gnd 54.00fF $ **FLOATING
C132 a_30384_802.n0 gnd 3.14fF $ **FLOATING
C133 a_38070_8852.n0 gnd 3.65fF $ **FLOATING
C134 a_50511_16072.n0 gnd 2.15fF $ **FLOATING
C135 a_28790_25040.n0 gnd 3.75fF $ **FLOATING
C136 a_32948_24994.n0 gnd 3.11fF $ **FLOATING
C137 a_23308_802.n0 gnd 3.31fF $ **FLOATING
C138 a_24410_25128.n0 gnd 3.81fF $ **FLOATING
C139 a_77254_23336.t2 gnd 36.73fF
C140 a_77254_23336.t4 gnd 56.94fF
C141 a_77254_23336.n0 gnd 60.94fF $ **FLOATING
C142 a_77254_23336.t3 gnd 44.97fF
C143 a_77254_23336.t1 gnd 65.92fF
C144 a_77254_23336.n1 gnd 94.34fF $ **FLOATING
C145 a_77254_23336.n2 gnd 94.36fF $ **FLOATING
C146 a_77254_23336.t0 gnd 38.38fF
C147 a_77254_23336.t5 gnd 41.73fF
C148 a_77254_23336.n3 gnd 14.94fF $ **FLOATING
C149 a_77254_23336.t6 gnd 3.54fF
C150 a_77280_24640.t2 gnd 28.50fF $ **FLOATING
C151 a_77280_24640.t4 gnd 36.40fF $ **FLOATING
C152 a_77280_24640.n0 gnd 62.35fF $ **FLOATING
C153 a_77280_24640.t1 gnd 36.30fF $ **FLOATING
C154 a_77280_24640.t3 gnd 44.53fF $ **FLOATING
C155 a_77280_24640.n1 gnd 24.73fF $ **FLOATING
C156 a_77280_24640.n2 gnd 126.44fF $ **FLOATING
C157 a_77280_24640.t0 gnd 2.47fF
C158 a_14910_6932.n0 gnd 3.12fF $ **FLOATING
C159 a_14832_12082.n0 gnd 3.86fF $ **FLOATING
C160 a_51138_19904.n0 gnd 2.56fF $ **FLOATING
C161 a_27762_11446.n0 gnd 4.89fF $ **FLOATING
C162 a_27762_11446.t47 gnd 9.88fF $ **FLOATING
C163 a_27762_11446.t21 gnd 9.88fF $ **FLOATING
C164 a_27762_11446.t11 gnd 7.39fF $ **FLOATING
C165 a_27762_11446.n3 gnd 12.90fF $ **FLOATING
C166 a_27762_11446.n4 gnd 4.16fF $ **FLOATING
C167 Fvco_By4_QPH_bar.n2 gnd 23.88fF $ **FLOATING
C168 Fvco_By4_QPH_bar.n4 gnd 3.41fF $ **FLOATING
C169 Fvco_By4_QPH_bar.n5 gnd 3.08fF $ **FLOATING
C170 Fvco_By4_QPH_bar.n7 gnd 6.96fF $ **FLOATING
C171 a_50583_13108.n0 gnd 8.05fF $ **FLOATING
C172 a_51516_3690.n1 gnd 3.35fF $ **FLOATING
C173 a_51516_3690.n2 gnd 3.11fF $ **FLOATING
C174 a_49916_3664.t1 gnd 4.56fF $ **FLOATING
C175 a_49858_3690.n0 gnd 4.03fF $ **FLOATING
C176 a_49858_3690.t5 gnd 2.40fF $ **FLOATING
C177 a_49858_3690.t7 gnd 2.45fF $ **FLOATING
C178 a_49858_3690.t8 gnd 2.24fF $ **FLOATING
C179 a_22429_17162.n0 gnd 3.53fF $ **FLOATING
C180 a_22429_17162.t34 gnd 46.82fF $ **FLOATING
C181 a_22429_17162.t29 gnd 10.84fF $ **FLOATING
C182 a_22429_17162.n1 gnd 7.36fF $ **FLOATING
C183 a_22429_17162.n3 gnd 4.66fF $ **FLOATING
C184 a_23436_16644.n0 gnd 4.67fF $ **FLOATING
C185 a_23436_16644.t60 gnd 10.21fF $ **FLOATING
C186 a_23436_16644.t12 gnd 8.90fF $ **FLOATING
C187 a_23436_16644.t46 gnd 6.39fF $ **FLOATING
C188 a_23436_16644.n3 gnd 3.27fF $ **FLOATING
C189 a_56334_20860.n0 gnd 2.57fF $ **FLOATING
C190 a_52052_20860.t18 gnd 3.50fF
C191 a_54432_7362.t1 gnd 3.00fF
C192 vbiasob.n2 gnd 6.14fF $ **FLOATING
C193 vbiasob.n3 gnd 5.05fF $ **FLOATING
C194 a_14266_8900.n0 gnd 4.92fF $ **FLOATING
C195 a_14266_8900.t54 gnd 9.27fF $ **FLOATING
C196 a_14266_8900.t47 gnd 9.98fF $ **FLOATING
C197 a_14266_8900.t16 gnd 12.27fF $ **FLOATING
C198 a_14266_8900.n4 gnd 10.34fF $ **FLOATING
C199 a_17685_3840.t18 gnd 2.78fF $ **FLOATING
C200 a_17685_3840.t59 gnd 2.78fF $ **FLOATING
C201 a_17685_3840.t54 gnd 2.78fF $ **FLOATING
C202 a_17685_3840.t56 gnd 2.78fF $ **FLOATING
C203 a_17685_3840.t49 gnd 2.78fF $ **FLOATING
C204 a_17685_3840.t44 gnd 2.78fF $ **FLOATING
C205 a_17685_3840.t16 gnd 2.78fF $ **FLOATING
C206 a_17685_3840.t60 gnd 2.78fF $ **FLOATING
C207 a_17685_3840.t52 gnd 2.78fF $ **FLOATING
C208 a_17685_3840.t47 gnd 2.78fF $ **FLOATING
C209 a_17685_3840.t39 gnd 6.44fF $ **FLOATING
C210 a_17685_3840.n1 gnd 11.36fF $ **FLOATING
C211 a_17685_3840.n2 gnd 7.40fF $ **FLOATING
C212 a_17685_3840.n3 gnd 7.40fF $ **FLOATING
C213 a_17685_3840.n4 gnd 7.40fF $ **FLOATING
C214 a_17685_3840.n5 gnd 7.40fF $ **FLOATING
C215 a_17685_3840.n6 gnd 7.40fF $ **FLOATING
C216 a_17685_3840.n7 gnd 7.40fF $ **FLOATING
C217 a_17685_3840.n8 gnd 7.40fF $ **FLOATING
C218 a_17685_3840.n9 gnd 7.40fF $ **FLOATING
C219 a_17685_3840.n10 gnd 6.25fF $ **FLOATING
C220 a_17685_3840.t50 gnd 3.74fF $ **FLOATING
C221 a_17685_3840.n11 gnd 7.66fF $ **FLOATING
C222 a_17685_3840.t42 gnd 2.78fF $ **FLOATING
C223 a_17685_3840.t34 gnd 2.78fF $ **FLOATING
C224 a_17685_3840.t27 gnd 2.78fF $ **FLOATING
C225 a_17685_3840.t29 gnd 2.78fF $ **FLOATING
C226 a_17685_3840.t20 gnd 2.78fF $ **FLOATING
C227 a_17685_3840.t14 gnd 2.78fF $ **FLOATING
C228 a_17685_3840.t57 gnd 2.78fF $ **FLOATING
C229 a_17685_3840.t51 gnd 2.78fF $ **FLOATING
C230 a_17685_3840.t45 gnd 2.78fF $ **FLOATING
C231 a_17685_3840.t38 gnd 2.78fF $ **FLOATING
C232 a_17685_3840.t31 gnd 6.44fF $ **FLOATING
C233 a_17685_3840.n12 gnd 11.34fF $ **FLOATING
C234 a_17685_3840.n13 gnd 7.39fF $ **FLOATING
C235 a_17685_3840.n14 gnd 7.39fF $ **FLOATING
C236 a_17685_3840.n15 gnd 7.39fF $ **FLOATING
C237 a_17685_3840.n16 gnd 7.39fF $ **FLOATING
C238 a_17685_3840.n17 gnd 7.39fF $ **FLOATING
C239 a_17685_3840.n18 gnd 7.39fF $ **FLOATING
C240 a_17685_3840.n19 gnd 7.39fF $ **FLOATING
C241 a_17685_3840.n20 gnd 7.39fF $ **FLOATING
C242 a_17685_3840.n21 gnd 6.25fF $ **FLOATING
C243 a_17685_3840.t23 gnd 3.74fF $ **FLOATING
C244 a_17685_3840.n22 gnd 5.61fF $ **FLOATING
C245 a_17685_3840.n23 gnd 6.37fF $ **FLOATING
C246 a_17685_3840.n24 gnd 3.21fF $ **FLOATING
C247 a_17685_3840.n27 gnd 2.54fF $ **FLOATING
C248 a_17685_3840.t43 gnd 2.78fF $ **FLOATING
C249 a_17685_3840.t37 gnd 2.78fF $ **FLOATING
C250 a_17685_3840.t40 gnd 2.78fF $ **FLOATING
C251 a_17685_3840.t32 gnd 2.78fF $ **FLOATING
C252 a_17685_3840.t25 gnd 2.78fF $ **FLOATING
C253 a_17685_3840.t24 gnd 2.78fF $ **FLOATING
C254 a_17685_3840.t17 gnd 2.78fF $ **FLOATING
C255 a_17685_3840.t58 gnd 2.78fF $ **FLOATING
C256 a_17685_3840.t53 gnd 2.78fF $ **FLOATING
C257 a_17685_3840.t46 gnd 6.44fF $ **FLOATING
C258 a_17685_3840.n32 gnd 11.32fF $ **FLOATING
C259 a_17685_3840.n33 gnd 7.38fF $ **FLOATING
C260 a_17685_3840.n34 gnd 7.38fF $ **FLOATING
C261 a_17685_3840.n35 gnd 7.38fF $ **FLOATING
C262 a_17685_3840.n36 gnd 7.38fF $ **FLOATING
C263 a_17685_3840.n37 gnd 7.38fF $ **FLOATING
C264 a_17685_3840.n38 gnd 7.38fF $ **FLOATING
C265 a_17685_3840.n39 gnd 7.38fF $ **FLOATING
C266 a_17685_3840.n40 gnd 7.38fF $ **FLOATING
C267 a_17685_3840.t48 gnd 2.78fF $ **FLOATING
C268 a_17685_3840.n41 gnd 6.22fF $ **FLOATING
C269 a_17685_3840.t35 gnd 3.75fF $ **FLOATING
C270 a_17685_3840.n42 gnd 7.71fF $ **FLOATING
C271 a_17685_3840.t41 gnd 2.78fF $ **FLOATING
C272 a_17685_3840.t33 gnd 2.78fF $ **FLOATING
C273 a_17685_3840.t26 gnd 2.78fF $ **FLOATING
C274 a_17685_3840.t28 gnd 2.78fF $ **FLOATING
C275 a_17685_3840.t19 gnd 2.78fF $ **FLOATING
C276 a_17685_3840.t13 gnd 2.78fF $ **FLOATING
C277 a_17685_3840.t36 gnd 2.78fF $ **FLOATING
C278 a_17685_3840.t30 gnd 2.78fF $ **FLOATING
C279 a_17685_3840.t21 gnd 2.78fF $ **FLOATING
C280 a_17685_3840.t15 gnd 2.78fF $ **FLOATING
C281 a_17685_3840.t55 gnd 6.44fF $ **FLOATING
C282 a_17685_3840.n43 gnd 11.37fF $ **FLOATING
C283 a_17685_3840.n44 gnd 7.41fF $ **FLOATING
C284 a_17685_3840.n45 gnd 7.41fF $ **FLOATING
C285 a_17685_3840.n46 gnd 7.41fF $ **FLOATING
C286 a_17685_3840.n47 gnd 7.41fF $ **FLOATING
C287 a_17685_3840.n48 gnd 7.41fF $ **FLOATING
C288 a_17685_3840.n49 gnd 7.41fF $ **FLOATING
C289 a_17685_3840.n50 gnd 7.41fF $ **FLOATING
C290 a_17685_3840.n51 gnd 7.41fF $ **FLOATING
C291 a_17685_3840.n52 gnd 6.26fF $ **FLOATING
C292 a_17685_3840.t22 gnd 3.74fF $ **FLOATING
C293 a_17685_3840.n53 gnd 5.43fF $ **FLOATING
C294 a_17685_3840.n54 gnd 6.25fF $ **FLOATING
C295 a_17685_3840.n55 gnd 3.40fF $ **FLOATING
C296 a_17685_3840.n60 gnd 2.24fF $ **FLOATING
C297 a_25099_11445.n0 gnd 4.85fF $ **FLOATING
C298 a_25099_11445.t40 gnd 9.08fF $ **FLOATING
C299 a_25099_11445.t15 gnd 10.03fF $ **FLOATING
C300 a_25099_11445.n3 gnd 2.56fF $ **FLOATING
C301 a_25099_11445.t53 gnd 8.63fF $ **FLOATING
C302 a_25099_11445.n4 gnd 7.06fF $ **FLOATING
C303 a_33804_31120.n6 gnd 33.76fF $ **FLOATING
C304 a_33804_31120.t4 gnd 5.96fF
C305 a_26036_4988.n0 gnd 9.29fF $ **FLOATING
C306 a_26036_4988.n1 gnd 4.19fF $ **FLOATING
C307 a_26036_4988.t20 gnd 9.20fF $ **FLOATING
C308 a_26036_4988.t44 gnd 6.43fF $ **FLOATING
C309 a_26036_4988.t16 gnd 5.98fF $ **FLOATING
C310 a_33900_31430.n16 gnd 43.12fF $ **FLOATING
C311 Fvco_By4_QPH.n0 gnd 11.17fF $ **FLOATING
C312 Fvco_By4_QPH.n7 gnd 2.17fF $ **FLOATING
C313 Fvco_By4_QPH.n8 gnd 2.14fF $ **FLOATING
C314 Fvco_By4_QPH.n9 gnd 4.51fF $ **FLOATING
C315 Fvco_By4_QPH.n11 gnd 4.92fF $ **FLOATING
C316 a_14188_14050.n0 gnd 9.38fF $ **FLOATING
C317 a_14188_14050.t39 gnd 4.60fF $ **FLOATING
C318 a_14188_14050.t31 gnd 20.11fF $ **FLOATING
C319 a_14188_14050.n3 gnd 3.53fF $ **FLOATING
C320 a_14188_14050.t12 gnd 10.19fF $ **FLOATING
C321 a_14188_14050.n4 gnd 10.20fF $ **FLOATING
C322 vinit.t40 gnd 14.88fF $ **FLOATING
C323 vinit.n18 gnd 210.62fF $ **FLOATING
C324 vinit.n28 gnd 2.88fF $ **FLOATING
C325 vinit.n29 gnd 2.86fF $ **FLOATING
C326 vbiasr.t40 gnd 28.85fF
C327 vbiasr.n16 gnd 119.71fF $ **FLOATING
C328 vbiasr.n27 gnd 4.28fF $ **FLOATING
C329 vbiasr.n28 gnd 4.24fF $ **FLOATING
C330 vbiasr.n39 gnd 3.21fF $ **FLOATING
C331 a_26690_784.n0 gnd 3.33fF $ **FLOATING
C332 a_23414_5032.n0 gnd 7.44fF $ **FLOATING
C333 a_23414_5032.t14 gnd 13.39fF $ **FLOATING
C334 a_23414_5032.n4 gnd 2.40fF $ **FLOATING
C335 a_23414_5032.t2 gnd 6.75fF $ **FLOATING
C336 a_23414_5032.n5 gnd 5.65fF $ **FLOATING
C337 a_26368_16652.n0 gnd 4.22fF $ **FLOATING
C338 a_26368_16652.t52 gnd 11.97fF $ **FLOATING
C339 a_26368_16652.t39 gnd 9.05fF $ **FLOATING
C340 a_26368_16652.t24 gnd 6.04fF $ **FLOATING
C341 a_26368_16652.n3 gnd 4.14fF $ **FLOATING
