* NGSPICE file created from a2.ext - technology: sky130A

X0 vdd a_34044_31208.t4 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1 vdd a_34044_31208.t5 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X2 Fvco_By4_QPH_bar.t1 a_66167_26022.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X3 a_28994_17218.t6 a_26368_16652.t2 a_28736_17218.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X4 a_26690_784.t1 a_23414_5032.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X5 vdd a_1026_45630.t4 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X6 vdd Vso1b.t2 a_4226_11420.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X7 a_28220_17218.t13 a_26368_16652.t3 a_27962_17218.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8 vdd a_34044_31208.t6 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X9 a_29510_17218.t6 a_26368_16652.t4 a_29252_17218.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X10 a_50320_14126.t2 Fvco_By4_QPH.t2 a_55602_11692.t5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_49874_4150.t0 a_49874_4150.t0 a_54950_4814.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.28e+06u l=8e+06u
X12 a_22629_5596.t6 a_14188_14050.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X13 a_23403_5596.t13 a_14188_14050.t3 a_23145_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X14 vdd a_1026_45630.t5 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X15 a_29510_17218.t5 a_26368_16652.t5 a_29252_17218.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X16 a_54950_4814.t0 a_49874_4150.t0 a_53292_4814.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.28e+06u l=8e+06u
X17 a_22887_5596.t6 a_14188_14050.t4 a_22629_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X18 a_28994_5597.t6 a_26036_4988.t2 a_28736_5597.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X19 a_1026_45630.t3 CLK_BY_4_IPH.t1 vctrl.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_26847_11500.t6 a_25099_11445.t2 a_26589_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X21 vdd a_66167_26022.t4 a_66154_26414.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X22 vdd a_1026_45630.t6 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X23 a_24177_5596.t12 a_14188_14050.t5 a_23919_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X24 vdd a_34044_31208.t7 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X25 gnd a_17685_3840.t17 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X26 a_22629_11500.t6 a_14266_8900.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X27 gnd a_17685_3840.t18 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X28 vdd a_34044_31208.t8 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X29 a_66357_25280.t0 RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X30 vdd a_34044_31208.t9 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X31 vdd a_63529_26290.t4 a_63419_26414.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X32 a_28736_5597.t8 a_26036_4988.t3 a_28478_5597.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X33 a_26847_11500.t5 a_25099_11445.t3 a_26589_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X34 a_29510_5597.t13 a_26036_4988.t4 a_29252_5597.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X35 vdd a_1026_45630.t7 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X36 gnd Vso3b.t2 a_8744_13422.t1 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X37 gnd a_17685_3840.t19 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X38 vdd a_1026_45630.t8 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X39 vdd a_1026_45630.t9 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X40 gnd Vso5b.t2 a_8748_12270.t1 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X41 a_26847_11500.t4 a_25099_11445.t4 a_26589_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X42 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X43 a_23919_5596.t4 a_14188_14050.t6 a_23661_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X44 a_28994_5597.t5 a_26036_4988.t5 a_28736_5597.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X45 vdd a_34044_31208.t10 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X46 vdd a_1026_45630.t10 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X47 a_52052_20860.t0 a_56334_20860.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X48 vdd a_34044_31208.t11 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X49 a_26847_11500.t3 a_25099_11445.t5 a_26589_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X50 a_23156_5032.t6 a_14188_14050.t7 a_24177_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X51 a_28736_17218.t2 a_26368_16652.t6 a_28478_17218.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X52 vdd a_34044_31208.t12 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X53 a_65546_25646.t0 RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X54 a_25299_17217.t6 a_23436_16644.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X55 vdd a_1026_45630.t11 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X56 vdd a_34044_31208.t13 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X57 vdd a_1026_45630.t12 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X58 a_26847_17217.t9 a_23436_16644.t3 a_26589_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X59 a_28736_17218.t13 a_26368_16652.t7 a_28478_17218.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X60 a_51276_14152.t3 Fvco_By4_QPH.t3 a_51636_13108.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 gnd a_17685_3840.t20 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X62 a_25815_5596.t8 a_23414_5032.t3 a_25557_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X63 vdd a_34044_31208.t14 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X64 vdd a_1026_45630.t13 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X65 a_63311_26048.t0 a_62795_26048.t2 a_63216_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X66 a_23145_5596.t11 a_14188_14050.t8 a_22887_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X67 a_26331_11500.t6 a_25099_11445.t6 a_26073_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X68 a_28478_5597.t1 a_26036_4988.t6 a_28220_5597.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X69 a_29252_5597.t12 a_26036_4988.t7 a_28994_5597.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X70 vdd a_34044_31208.t15 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X71 vdd a_34044_31208.t16 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X72 vdd CLK_IN.t2 a_4288_11534.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X73 a_25778_4988.t7 a_23414_5032.t4 a_26847_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X74 vdd a_1026_45630.t14 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X75 vdd a_34044_31208.t17 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X76 a_26331_11500.t5 a_25099_11445.t7 a_26073_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X77 gnd a_17685_3840.t21 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X78 a_23145_17217.t6 Fvco.t2 a_22887_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X79 vdd a_1026_45630.t15 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X80 vdd a_34044_31208.t18 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X81 vdd a_1026_45630.t16 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X82 vdd a_34044_31208.t19 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X83 a_28220_17218.t12 a_26368_16652.t8 a_27962_17218.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X84 a_23145_17217.t5 Fvco.t3 a_22887_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X85 a_52052_20860.t5 a_51636_13108.t5 a_56602_11692.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X86 a_56602_11692.t13 vbiasob.t3 a_56272_15934.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X87 a_27962_5597.t6 a_26036_4988.t8 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X88 vdd a_34044_31208.t20 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X89 vbiasbuffer.t2 a_49874_4150.t0 a_54966_2992.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=8e+06u
X90 vdd a_1026_45630.t17 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X91 vdd a_1026_45630.t18 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X92 a_26331_17217.t6 a_23436_16644.t4 a_26073_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X93 a_28220_17218.t11 a_26368_16652.t9 a_27962_17218.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X94 vbiasob.t2 a_57726_5786.t5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.40205e+11p ps=1.78513e+06u w=1.02e+06u l=1e+06u
X95 a_25557_11500.t12 a_25099_11445.t8 a_25299_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X96 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X97 a_25557_5596.t10 a_23414_5032.t5 a_25299_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X98 a_22887_5596.t5 a_14188_14050.t9 a_22629_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X99 a_23661_5596.t6 a_14188_14050.t10 a_23403_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X100 vdd a_34044_31208.t21 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X101 vdd a_1026_45630.t19 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X102 a_26847_5596.t0 a_23414_5032.t6 a_26589_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X103 vdd a_34044_31208.t22 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X104 a_28578_5014.t7 a_26036_4988.t9 a_29510_5597.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X105 vdd a_1026_45630.t20 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X106 gnd a_17685_3840.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X107 a_28220_5597.t13 a_26036_4988.t10 a_27962_5597.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X108 vdd a_34044_31208.t23 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X109 a_24177_11500.t6 a_14266_8900.t3 a_23919_11500.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X110 a_50583_13108.t1 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X111 a_25557_11500.t11 a_25099_11445.t9 a_25299_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X112 a_52052_20860.t17 a_51041_13108.t5 a_55602_11692.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X113 a_23403_5596.t12 a_14188_14050.t11 a_23145_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X114 vdd a_1026_45630.t21 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X115 a_29252_11501.t13 a_27762_11446.t2 a_28994_11501.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X116 a_25557_11500.t10 a_25099_11445.t10 a_25299_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X117 a_25299_5596.t6 a_23414_5032.t7 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X118 vdd a_34044_31208.t24 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X119 a_49932_4124.t1 a_49932_4124.t0 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=2e+07u
X120 a_28994_5597.t4 a_26036_4988.t11 a_28736_5597.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X121 vdd a_1026_45630.t22 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X122 vdd a_1026_45630.t23 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X123 a_25557_11500.t9 a_25099_11445.t11 a_25299_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X124 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X125 a_65438_25280.t2 a_65088_25280.t2 a_65343_25280.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X126 a_66346_26048.t0 RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X127 a_26589_5596.t0 a_23414_5032.t8 a_26331_5596.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X128 vdd a_34044_31208.t25 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X129 a_65656_25522.t1 a_65438_25280.t4 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.27414e+11p ps=920615u w=840000u l=150000u
X130 a_24177_11500.t5 a_14266_8900.t4 a_23919_11500.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X131 a_44752_16348.t2 a_51138_19904.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X132 a_25557_17217.t7 a_23436_16644.t5 a_25299_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X133 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X134 vdd a_1026_45630.t24 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X135 vdd a_34044_31208.t26 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X136 a_24177_11500.t4 a_14266_8900.t5 a_23919_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X137 a_27962_11501.t6 a_27762_11446.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X138 vdd a_1026_45630.t25 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X139 a_14832_12082.t1 a_14188_14050.t12 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X140 a_29252_11501.t12 a_27762_11446.t4 a_28994_11501.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X141 a_56602_11692.t11 a_51636_13108.t6 a_52052_20860.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X142 a_29510_5597.t12 a_26036_4988.t12 a_29252_5597.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X143 a_24177_11500.t3 a_14266_8900.t6 a_23919_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X144 vdd a_34044_31208.t27 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X145 zz.t0 CLK_BY_4_IPH_BAR.t0 a_34044_31208.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X146 a_66003_25280.t1 a_64922_25280.t2 a_65656_25522.t3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X147 a_29252_11501.t11 a_27762_11446.t5 a_28994_11501.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X148 vdd a_56334_19906.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X149 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X150 a_26073_5596.t13 a_23414_5032.t9 a_25815_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X151 vdd a_1026_45630.t26 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X152 vdd a_34044_31208.t28 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X153 a_24177_17217.t10 Fvco.t4 a_23919_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X154 a_29252_11501.t10 a_27762_11446.t6 a_28994_11501.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X155 a_26847_17217.t8 a_23436_16644.t6 a_26589_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X156 a_23160_10936.t7 a_14266_8900.t7 a_24177_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X157 vdd a_34044_31208.t29 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X158 gnd Vso7b.t2 a_8748_11114.t1 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X159 a_29252_17218.t6 a_26368_16652.t10 a_28994_17218.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X160 a_23661_11500.t13 a_14266_8900.t8 a_23403_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X161 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X162 a_26847_17217.t7 a_23436_16644.t7 a_26589_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X163 vdd a_34044_31208.t30 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X164 a_23661_11500.t12 a_14266_8900.t9 a_23403_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X165 a_25815_5596.t7 a_23414_5032.t10 a_25557_5596.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X166 a_23919_11500.t11 a_14266_8900.t10 a_23661_11500.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X167 a_26331_5596.t9 a_23414_5032.t11 a_26073_5596.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X168 a_55602_11692.t12 a_51041_13108.t6 a_52052_20860.t18 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X169 a_42574_15624.t2 Fvco_By4_QPH_bar.t2 a_42550_16062.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X170 a_29252_5597.t11 a_26036_4988.t13 a_28994_5597.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X171 a_53308_3580.t0 a_49874_4150.t0 vbiasr.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.83e+06u l=8e+06u
X172 vdd a_1026_45630.t27 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X173 a_23661_17217.t13 Fvco.t5 a_23403_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X174 vdd a_34044_31208.t31 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X175 a_26331_17217.t5 a_23436_16644.t8 a_26073_17217.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X176 a_22887_11500.t6 a_14266_8900.t11 a_22629_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X177 CLK_BY_4_IPH_BAR a_66742_25280.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X178 a_28438_10874.t7 a_27762_11446.t7 a_29510_11501.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X179 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X180 vdd a_34044_31208.t32 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X181 gnd a_17685_3840.t23 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X182 a_26331_17217.t4 a_23436_16644.t9 a_26073_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X183 a_23919_11500.t13 a_14266_8900.t12 a_23661_11500.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X184 gnd a_17685_3840.t24 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X185 vdd a_1026_45630.t28 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X186 a_28438_10874.t6 a_27762_11446.t8 a_29510_11501.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X187 a_25557_5596.t9 a_23414_5032.t12 a_25299_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X188 a_23919_11500.t12 a_14266_8900.t13 a_23661_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X189 vdd a_34044_31208.t33 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X190 a_65438_25280.t3 a_64922_25280.t3 a_65343_25280.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X191 a_23919_11500.t8 a_14266_8900.t14 a_23661_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X192 vdd a_34044_31208.t34 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X193 a_63573_26048.t1 a_63529_26290.t5 a_63407_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X194 gnd a_17685_3840.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X195 a_22887_11500.t5 a_14266_8900.t15 a_22629_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X196 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X197 vdd a_34044_31208.t35 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X198 vdd a_34044_31208.t36 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X199 a_14910_6932.t1 a_14266_8900.t16 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X200 vdd a_1026_45630.t29 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X201 a_28622_16652.t6 a_26368_16652.t11 a_29510_17218.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X202 vdd a_1026_45630.t30 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X203 gnd Vso4b.t2 a_8740_12844.t0 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X204 a_4314_11564.t0 a_4288_11534.t3 a_4314_11468.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X205 a_23919_17217.t6 Fvco.t6 a_23661_17217.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X206 a_22887_11500.t4 a_14266_8900.t17 a_22629_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X207 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X208 vdd a_34044_31208.t37 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X209 gnd a_17685_3840.t26 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X210 gnd a_17685_3840.t27 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X211 vdd a_1026_45630.t31 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X212 vdd a_4288_11918.t3 vout.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X213 a_23403_11500.t7 a_14266_8900.t18 a_23145_11500.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X214 a_22887_11500.t3 a_14266_8900.t19 a_22629_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X215 CLK_BY_2_BAR.t0 a_64615_26048.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X216 vdd a_1026_45630.t32 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X217 a_23403_11500.t13 a_14266_8900.t20 a_23145_11500.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X218 a_26016_10878.t6 a_25099_11445.t12 a_26847_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X219 a_25299_5596.t5 a_23414_5032.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X220 vdd a_34044_31208.t38 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X221 a_22887_17217.t2 Fvco.t7 a_22629_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X222 a_64725_25280.t3 CLK_BY_2_BAR.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X223 a_28622_16652.t5 a_26368_16652.t12 a_29510_17218.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X224 vdd a_34044_31208.t39 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X225 a_25557_17217.t6 a_23436_16644.t10 a_25299_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X226 vdd a_1026_45630.t33 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X227 gnd a_17685_3840.t28 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X228 a_25557_17217.t5 a_23436_16644.t11 a_25299_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X229 a_26073_11500.t5 a_25099_11445.t13 a_25815_11500.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X230 gnd a_57726_5786.t3 a_57726_5786.t4 gnd sky130_fd_pr__nfet_01v8 ad=7.06485e+11p pd=5.25039e+06u as=0p ps=0u w=3e+06u l=1e+06u
X231 vdd a_1026_45630.t34 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X232 a_23403_17217.t13 Fvco.t8 a_23145_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X233 vdd a_1026_45630.t35 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X234 vdd a_34044_31208.t40 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X235 a_22629_11500.t5 a_14266_8900.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X236 vdd a_1026_45630.t36 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X237 a_49932_4124.t2 a_49874_4150.t0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.01433e+11p ps=2.24017e+06u w=1.28e+06u l=8e+06u
X238 vdd a_34044_31208.t41 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X239 a_24177_17217.t9 Fvco.t9 a_23919_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X240 vdd a_1026_45630.t37 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X241 vdd a_1026_45630.t38 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X242 a_24177_17217.t8 Fvco.t10 a_23919_17217.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X243 vdd a_34044_31208.t42 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X244 gnd RESET a_63573_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X245 a_29252_17218.t5 a_26368_16652.t13 a_28994_17218.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X246 vbiasob.t1 vbiasob.t0 a_54448_7822.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X247 vdd a_34044_31208.t43 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X248 Vso1b.t1 a_24410_25128.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X249 a_28478_11501.t12 a_27762_11446.t9 a_28220_11501.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X250 a_29252_17218.t4 a_26368_16652.t14 a_28994_17218.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X251 a_22629_11500.t4 a_14266_8900.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X252 a_23308_802.t0 Fvco.t11 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X253 vdd a_1026_45630.t39 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X254 vdd a_1026_45630.t40 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X255 vdd a_34044_31208.t44 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X256 a_26368_16652.t1 a_23436_16644.t12 a_26110_16652.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X257 a_28478_11501.t11 a_27762_11446.t10 a_28220_11501.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X258 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.35495e+11p pd=1.75013e+06u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X259 a_24177_5596.t11 a_14188_14050.t13 a_23919_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X260 vdd a_1026_45630.t41 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X261 a_22629_11500.t3 a_14266_8900.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X262 a_22629_11500.t2 a_14266_8900.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X263 vdd a_34044_31208.t45 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X264 a_23661_17217.t12 Fvco.t12 a_23403_17217.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X265 gnd Vso1b.t3 a_8744_9386.t0 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X266 a_28478_17218.t13 a_26368_16652.t15 a_28220_17218.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X267 vdd a_34044_31208.t46 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X268 vdd a_1026_45630.t42 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X269 a_22629_17217.t6 Fvco.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X270 a_23661_17217.t11 Fvco.t14 a_23403_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X271 a_26036_4988.t1 a_23414_5032.t14 a_17685_3840.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X272 vdd a_34044_31208.t47 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X273 vdd a_4226_11420.t3 vout.t6 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X274 vdd a_1026_45630.t43 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X275 gnd a_64725_25280.t4 a_64922_25280.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X276 vdd a_34044_31208.t48 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X277 vdd a_34044_31208.t49 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X278 vdd a_4226_12188.t3 vout.t4 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X279 a_25815_11500.t13 a_25099_11445.t14 a_25557_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X280 vdd a_34044_31208.t50 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X281 vdd a_34044_31208.t51 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X282 a_32948_24994.t1 a_27762_11446.t11 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X283 Vso2b.t0 a_28790_25040.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X284 a_28478_17218.t12 a_26368_16652.t16 a_28220_17218.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X285 vdd a_1026_45630.t44 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X286 a_28622_16652.t4 a_26368_16652.t17 a_29510_17218.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X287 a_23145_5596.t10 a_14188_14050.t14 a_22887_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X288 a_23919_17217.t5 Fvco.t15 a_23661_17217.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X289 vdd a_34044_31208.t52 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X290 gnd a_17685_3840.t29 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X291 a_28622_16652.t3 a_26368_16652.t18 a_29510_17218.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X292 vdd a_66167_26022.t5 a_66731_26048.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=9.70773e+10p pd=701421u as=0p ps=0u w=640000u l=150000u
X293 a_23919_17217.t11 Fvco.t16 a_23661_17217.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X294 a_14910_6932.t0 a_14266_8900.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X295 gnd a_17685_3840.t30 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X296 a_52052_20860.t1 a_51636_13108.t7 a_56602_11692.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X297 gnd a_17685_3840.t31 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X298 vdd a_34044_31208.t53 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X299 a_51276_14152.t9 a_51334_14126.t4 z.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X300 vdd a_65992_26048.t4 a_66167_26022.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X301 vdd Vso6b.t2 a_4226_11804.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X302 a_22887_17217.t8 Fvco.t17 a_22629_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X303 a_29510_11501.t13 a_27762_11446.t12 a_29252_11501.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X304 a_27962_5597.t5 a_26036_4988.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X305 vdd a_1026_45630.t45 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X306 vdd a_1026_45630.t46 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X307 a_22887_17217.t9 Fvco.t18 a_22629_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X308 a_51532_4150.t2 a_51532_4150.t1 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.51794e+11p ps=1.81931e+06u w=1.66e+06u l=4e+06u
X309 vdd a_1026_45630.t47 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X310 vdd a_65656_25522.t4 a_65546_25646.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X311 vdd CLK_BY_2_BAR.t3 a_64911_26048.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=9.70773e+10p pd=701421u as=0p ps=0u w=640000u l=150000u
X312 a_56602_11692.t9 a_51636_13108.t8 a_52052_20860.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X313 vdd a_50032_16080.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X314 vdd a_34044_31208.t54 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X315 a_23403_17217.t12 Fvco.t19 a_23145_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X316 a_50511_16072.t5 a_50320_14126.t4 a_50262_14152.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X317 a_22887_5596.t4 a_14188_14050.t15 a_22629_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X318 a_23661_5596.t5 a_14188_14050.t16 a_23403_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X319 vdd a_1026_45630.t48 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X320 a_64038_26414.t0 a_62961_26048.t2 a_63876_26048.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X321 a_23403_17217.t11 Fvco.t20 a_23145_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X322 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X323 vdd a_51138_19904.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X324 a_23919_5596.t3 a_14188_14050.t17 a_23661_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X325 z.t6 a_51334_14126.t5 a_51276_14152.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X326 vdd a_1026_45630.t49 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X327 a_52052_20860.t13 a_51041_13108.t7 a_55602_11692.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X328 a_50583_13108.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X329 vdd a_34044_31208.t55 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X330 vdd a_1026_45630.t50 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X331 vdd a_1026_45630.t51 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X332 a_65534_25280.t0 a_65088_25280.t3 a_65438_25280.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X333 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X334 a_27962_11501.t5 a_27762_11446.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X335 Vso4b.t0 a_38070_8852.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X336 a_52052_20224.t0 a_56272_15934.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X337 vdd a_34044_31208.t56 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X338 vdd a_34044_31208.t57 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X339 a_14266_8900.t1 a_25099_11445.t15 a_26016_10878.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X340 vdd a_1026_45630.t52 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X341 a_28994_5597.t3 a_26036_4988.t15 a_28736_5597.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X342 Vso5b.t0 a_14910_6932.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X343 a_26589_11500.t6 a_25099_11445.t16 a_26331_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X344 a_55602_11692.t8 a_51041_13108.t8 a_52052_20860.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X345 a_26589_11500.t5 a_25099_11445.t17 a_26331_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X346 a_24177_5596.t10 a_14188_14050.t18 a_23919_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X347 a_23919_5596.t6 a_14188_14050.t19 a_23661_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X348 vdd a_34044_31208.t58 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X349 vdd a_34044_31208.t59 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X350 vdd a_1026_45630.t53 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X351 vdd a_1026_45630.t54 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X352 Fvco_By4_QPH_bar.t0 a_66167_26022.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X353 a_23160_10936.t6 a_14266_8900.t26 a_24177_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X354 a_27962_11501.t4 a_27762_11446.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X355 a_64230_26048.t0 RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X356 a_56602_11692.t8 a_51636_13108.t9 a_52052_20860.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X357 a_27962_11501.t3 a_27762_11446.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X358 a_28478_17218.t11 a_26368_16652.t19 a_28220_17218.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X359 z.t5 a_51334_14126.t6 a_51276_14152.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X360 a_30384_802.t1 a_26036_4988.t16 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X361 vdd a_34044_31208.t60 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X362 a_4314_12044.t0 a_4226_11996.t3 a_4314_11948.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X363 a_26589_17217.t6 a_23436_16644.t13 a_26331_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X364 a_22629_17217.t5 Fvco.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X365 a_27962_11501.t2 a_27762_11446.t16 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X366 vdd a_34044_31208.t61 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X367 gnd CLK_BY_2_BAR.t4 a_64911_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X368 a_65656_25522.t0 a_65438_25280.t5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.50717e+11p ps=1.12008e+06u w=640000u l=150000u
X369 a_28478_17218.t10 a_26368_16652.t20 a_28220_17218.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X370 a_26073_5596.t12 a_23414_5032.t15 a_25815_5596.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X371 vdd a_1026_45630.t55 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X372 a_22629_17217.t4 Fvco.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X373 a_23145_11500.t13 a_14266_8900.t27 a_22887_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X374 a_23160_10936.t5 a_14266_8900.t28 a_24177_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X375 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X376 vdd a_34044_31208.t62 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X377 a_27962_17218.t6 a_26368_16652.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X378 a_51041_13108.t4 a_50511_16072.t8 a_50583_13108.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X379 vdd a_34044_31208.t63 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X380 a_66167_26022.t0 RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X381 a_23160_10936.t4 a_14266_8900.t29 a_24177_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X382 a_28220_11501.t12 a_27762_11446.t17 a_27962_11501.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X383 a_57726_5786.t0 a_51532_4150.t4 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.60895e+11p ps=1.88507e+06u w=1.72e+06u l=4e+06u
X384 a_28578_5014.t6 a_26036_4988.t17 a_29510_5597.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X385 vdd a_1026_45630.t56 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X386 a_23160_10936.t3 a_14266_8900.t30 a_24177_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X387 vdd a_34044_31208.t64 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X388 vdd a_34044_31208.t65 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X389 a_26847_17217.t6 a_23436_16644.t14 a_26589_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X390 vdd a_1026_45630.t57 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X391 a_63311_26048.t2 a_62961_26048.t3 a_63216_26048.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X392 a_55602_11692.t9 a_51041_13108.t9 a_52052_20860.t15 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X393 vdd a_34044_31208.t66 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X394 a_65088_25280.t1 a_64922_25280.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X395 vdd a_54410_8156.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X396 a_23403_5596.t11 a_14188_14050.t20 a_23145_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X397 vdd a_1026_45630.t58 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X398 vdd a_1026_45630.t59 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X399 a_23178_16644.t7 Fvco.t23 a_24177_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X400 CLK_IN.t1 a_23308_802.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X401 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X402 a_50128_8156.t1 a_54448_7822.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X403 vdd a_1026_45630.t60 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X404 a_65546_25646.t1 a_64922_25280.t5 a_65438_25280.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X405 gnd a_17685_3840.t32 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X406 a_53308_2992.t0 a_49874_4150.t0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.17918e+11p ps=2.36268e+06u w=1.35e+06u l=8e+06u
X407 gnd a_17685_3840.t33 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X408 vdd a_1026_45630.t61 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X409 a_28578_5014.t5 a_26036_4988.t18 a_29510_5597.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X410 vdd a_1026_45630.t62 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X411 gnd Vso2b.t2 a_8736_14034.t1 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X412 a_27962_5597.t4 a_26036_4988.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X413 vdd a_34044_31208.t67 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X414 vdd a_1026_45630.t63 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X415 vdd a_4226_11996.t4 vout.t3 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X416 vdd a_1026_45630.t64 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X417 vdd a_34044_31208.t68 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X418 vdd a_34044_31208.t69 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X419 gnd a_17685_3840.t34 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X420 Fvco.t0 a_26036_4988.t20 a_28578_5014.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X421 a_22629_5596.t5 a_14188_14050.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X422 a_26016_10878.t5 a_25099_11445.t18 a_26847_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X423 a_25299_11500.t6 a_25099_11445.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X424 a_23403_5596.t10 a_14188_14050.t22 a_23145_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X425 a_29510_5597.t11 a_26036_4988.t21 a_29252_5597.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X426 a_17685_3840.t11 vinit vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=1e+06u
X427 a_23661_5596.t4 a_14188_14050.t23 a_23403_5596.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X428 vdd a_63876_26048.t4 a_64051_26022.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X429 a_25299_11500.t5 a_25099_11445.t20 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X430 a_23919_5596.t5 a_14188_14050.t24 a_23661_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X431 vdd a_1026_45630.t65 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X432 vdd a_1026_45630.t66 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X433 vdd a_34044_31208.t70 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X434 gnd a_17685_3840.t35 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X435 vdd a_1026_45630.t67 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X436 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X437 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X438 a_26073_11500.t12 a_25099_11445.t21 a_25815_11500.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X439 a_65077_26048.t1 a_64911_26048.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.70773e+10p ps=701421u w=640000u l=150000u
X440 a_25299_17217.t5 a_23436_16644.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X441 Vso7b.t1 a_26690_784.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X442 a_30384_802.t0 a_26036_4988.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X443 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X444 vdd a_1026_45630.t68 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X445 a_26016_10878.t4 a_25099_11445.t22 a_26847_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X446 a_25815_5596.t6 a_23414_5032.t16 a_25557_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X447 a_28736_5597.t7 a_26036_4988.t23 a_28478_5597.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X448 vdd a_1026_45630.t69 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X449 a_26016_10878.t3 a_25099_11445.t23 a_26847_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X450 a_29510_5597.t10 a_26036_4988.t24 a_29252_5597.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X451 a_29252_5597.t10 a_26036_4988.t25 a_28994_5597.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X452 vdd a_34044_31208.t71 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X453 vdd a_1026_45630.t70 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X454 a_66112_25280.t0 a_64922_25280.t6 a_66003_25280.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X455 a_26016_10878.t2 a_25099_11445.t24 a_26847_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X456 gnd a_17685_3840.t36 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X457 a_26073_11500.t7 a_25099_11445.t25 a_25815_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X458 a_56602_11692.t0 Fvco_By4_QPH_bar.t3 a_50320_14126.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X459 a_23156_5032.t5 a_14188_14050.t25 a_24177_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X460 gnd a_17685_3840.t37 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X461 a_46856_21176.t1 a_51138_21494.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X462 gnd a_17685_3840.t38 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X463 vdd a_1026_45630.t71 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X464 vdd a_34044_31208.t72 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X465 a_26110_16652.t6 a_23436_16644.t16 a_26847_17217.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X466 a_25557_17217.t4 a_23436_16644.t17 a_25299_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X467 a_26073_11500.t9 a_25099_11445.t26 a_25815_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X468 a_65645_26290.t1 a_65427_26048.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.50717e+11p ps=1.12008e+06u w=640000u l=150000u
X469 a_26589_17217.t11 a_23436_16644.t18 a_26331_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X470 a_26073_11500.t8 a_25099_11445.t27 a_25815_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X471 a_26589_17217.t10 a_23436_16644.t19 a_26331_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X472 a_25815_5596.t5 a_23414_5032.t17 a_25557_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X473 vdd a_34044_31208.t73 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X474 a_27962_17218.t5 a_26368_16652.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X475 a_42574_15624.t6 vbiasot.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=4e+06u
X476 gnd a_56334_20860.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X477 a_26073_5596.t11 a_23414_5032.t18 a_25815_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X478 a_28478_5597.t0 a_26036_4988.t26 a_28220_5597.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X479 a_25557_5596.t12 a_23414_5032.t19 a_25299_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X480 vdd a_34044_31208.t74 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X481 gnd a_64051_26022.t3 a_64615_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X482 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X483 a_29252_5597.t9 a_26036_4988.t27 a_28994_5597.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X484 a_26073_17217.t1 a_23436_16644.t20 a_25815_17217.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X485 a_24177_17217.t7 Fvco.t24 a_23919_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X486 a_27962_17218.t4 a_26368_16652.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X487 a_25778_4988.t6 a_23414_5032.t20 a_26847_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X488 gnd a_17685_3840.t39 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X489 a_26331_11500.t4 a_25099_11445.t28 a_26073_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X490 vdd a_1026_45630.t72 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X491 vdd vinit a_17685_3840.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51683e+11p pd=1.09597e+06u as=0p ps=0u w=1e+06u l=1e+06u
X492 a_28578_5014.t4 a_26036_4988.t28 a_29510_5597.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X493 vdd a_34044_31208.t75 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X494 a_65077_26048.t0 a_64911_26048.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X495 vdd Vso3b.t3 a_4288_12110.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X496 vdd a_34044_31208.t76 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X497 vdd a_34044_31208.t77 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X498 vdd a_34044_31208.t78 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X499 vdd CLK_BY_2_BAR.t5 a_64725_25280.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=1.51683e+11p pd=1.09597e+06u as=0p ps=0u w=1e+06u l=150000u
X500 vdd Vso5b.t3 a_4288_11918.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X501 a_23178_16644.t6 Fvco.t25 a_24177_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X502 a_34044_31208.t2 CLK_BY_4_IPH.t2 zz.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X503 Vso3b.t0 a_32948_24994.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X504 a_25815_11500.t12 a_25099_11445.t29 a_25557_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X505 a_23403_5596.t9 a_14188_14050.t26 a_23145_5596.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X506 vdd a_34044_31208.t79 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X507 a_23178_16644.t5 Fvco.t26 a_24177_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X508 a_25557_5596.t11 a_23414_5032.t21 a_25299_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X509 vdd a_1026_45630.t73 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X510 vdd a_1026_45630.t74 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X511 a_23504_23306.t1 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X512 a_25299_5596.t4 a_23414_5032.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X513 vdd a_1026_45630.t75 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X514 zz.t1 CLK_BY_4_IPH_BAR.t1 a_1026_45630.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X515 a_51636_13108.t4 a_50511_16072.t9 a_46856_19268.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X516 a_26847_5596.t13 a_23414_5032.t23 a_26589_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X517 vdd a_1026_45630.t76 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X518 vdd a_34044_31208.t80 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X519 a_25815_11500.t11 a_25099_11445.t30 a_25557_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X520 bb.t3 Fvco_By4_QPH.t4 a_47968_16078.t3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X521 a_28220_5597.t12 a_26036_4988.t29 a_27962_5597.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X522 vdd a_34044_31208.t81 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X523 vdd Vso7b.t3 a_4226_11612.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X524 vdd a_1026_45630.t77 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X525 a_29510_11501.t12 a_27762_11446.t18 a_29252_11501.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X526 a_25815_11500.t10 a_25099_11445.t31 a_25557_11500.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X527 vdd a_1026_45630.t78 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X528 vdd a_34044_31208.t82 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X529 a_29510_5597.t9 a_26036_4988.t30 a_29252_5597.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X530 a_25815_11500.t9 a_25099_11445.t32 a_25557_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X531 a_47968_16078.t1 Fvco_By4_QPH_bar.t4 aa.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X532 a_25299_5596.t3 a_23414_5032.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X533 vdd a_1026_45630.t79 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X534 vdd a_1026_45630.t80 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X535 vdd a_34044_31208.t83 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X536 Vso3b.t1 a_32948_24994.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X537 vdd a_34044_31208.t84 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X538 vdd a_1026_45630.t81 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X539 vdd Vso7b.t4 a_4288_11726.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X540 a_25815_17217.t13 a_23436_16644.t21 a_25557_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X541 a_25299_17217.t4 a_23436_16644.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X542 a_26589_5596.t2 a_23414_5032.t25 a_26331_5596.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X543 vdd a_1026_45630.t82 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X544 a_23919_17217.t10 Fvco.t27 a_23661_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X545 a_1026_45630.t2 CLK_BY_4_IPH.t3 zz.t3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X546 a_25299_17217.t3 a_23436_16644.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X547 a_29510_11501.t11 a_27762_11446.t19 a_29252_11501.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X548 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X549 a_25815_5596.t4 a_23414_5032.t26 a_25557_5596.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X550 vdd a_34044_31208.t85 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X551 vdd a_1026_45630.t83 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X552 a_63407_26048.t1 a_62961_26048.t4 a_63311_26048.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X553 a_29510_11501.t10 a_27762_11446.t20 a_29252_11501.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X554 CLK_IN.t0 a_23308_802.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X555 vdd a_34044_31208.t86 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X556 vdd a_1026_45630.t84 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X557 a_66101_26048.t0 a_64911_26048.t4 a_65992_26048.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X558 a_25099_11445.t1 a_27762_11446.t21 a_28438_10874.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X559 a_28790_25040.t1 a_26368_16652.t24 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X560 a_22887_17217.t1 Fvco.t28 a_22629_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X561 a_29510_11501.t9 a_27762_11446.t22 a_29252_11501.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X562 a_29252_5597.t8 a_26036_4988.t31 a_28994_5597.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X563 vdd a_1026_45630.t85 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X564 a_65535_26414.t2 RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X565 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X566 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X567 vdd a_34044_31208.t87 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X568 vdd a_34044_31208.t88 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X569 a_26110_16652.t5 a_23436_16644.t24 a_26847_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X570 vdd a_34044_31208.t89 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X571 vdd a_1026_45630.t86 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X572 vdd a_1026_45630.t87 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X573 Vso5b.t1 a_14910_6932.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X574 a_23436_16644.t1 Fvco.t29 a_17685_3840.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X575 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X576 vbiasot.t2 vbiasot.t1 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=4e+06u
X577 vdd a_1026_45630.t88 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X578 a_29510_17218.t4 a_26368_16652.t25 a_29252_17218.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X579 Vso7b.t0 a_26690_784.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X580 vdd a_1026_45630.t89 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X581 a_26110_16652.t4 a_23436_16644.t25 a_26847_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X582 vdd a_34044_31208.t90 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X583 vdd a_1026_45630.t90 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X584 a_23661_11500.t11 a_14266_8900.t31 a_23403_11500.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X585 vdd a_1026_45630.t91 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X586 vdd a_1026_45630.t92 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X587 vdd a_1026_45630.t93 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X588 a_26073_17217.t4 a_23436_16644.t26 a_25815_17217.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X589 a_25557_5596.t8 a_23414_5032.t27 a_25299_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X590 vdd Vso8b.t2 a_4288_11534.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X591 a_26331_5596.t8 a_23414_5032.t28 a_26073_5596.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X592 gnd a_17685_3840.t40 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X593 a_26073_17217.t8 a_23436_16644.t27 a_25815_17217.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X594 gnd a_17685_3840.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X595 a_50262_14152.t2 Fvco_By4_QPH.t5 a_51041_13108.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X596 a_47968_16078.t5 a_42550_16062.t4 a_50511_16072.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X597 CLK_BY_2.t1 a_64051_26022.t4 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X598 a_23145_11500.t12 a_14266_8900.t32 a_22887_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X599 a_49874_4150.t1 a_51532_4150.t5 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.51794e+11p ps=1.81931e+06u w=1.66e+06u l=4e+06u
X600 vdd CLK_IN.t3 a_4226_11420.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X601 vdd a_34044_31208.t91 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X602 vdd a_1026_45630.t94 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X603 bb.t2 vbiasbuffer.t3 a_51826_16054.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X604 vdd a_1026_45630.t95 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X605 a_28220_11501.t11 a_27762_11446.t23 a_27962_11501.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X606 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X607 vdd a_34044_31208.t92 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X608 vdd a_34044_31208.t93 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X609 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.29693e+12p pd=2.45018e+07u as=3.29693e+12p ps=2.45018e+07u w=1.4e+07u l=1e+06u
X610 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X611 vdd a_34044_31208.t94 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X612 a_28438_10874.t5 a_27762_11446.t24 a_29510_11501.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X613 a_43010_16058.t3 Fvco_By4_QPH.t6 a_42574_15624.t4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X614 a_25299_5596.t2 a_23414_5032.t29 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X615 Fvco_By4_QPH.t0 a_66731_26048.t2 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X616 a_28994_11501.t9 a_27762_11446.t25 a_28736_11501.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X617 a_23145_11500.t11 a_14266_8900.t33 a_22887_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X618 a_22629_17217.t3 Fvco.t30 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X619 a_28994_11501.t12 a_27762_11446.t26 a_28736_11501.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X620 a_23145_11500.t10 a_14266_8900.t34 a_22887_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X621 a_28220_11501.t10 a_27762_11446.t27 a_27962_11501.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X622 vdd a_1026_45630.t96 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X623 a_23145_11500.t9 a_14266_8900.t35 a_22887_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X624 a_50511_16072.t4 a_50320_14126.t5 a_50262_14152.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X625 vdd a_34044_31208.t95 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X626 a_66165_25646.t0 a_65088_25280.t4 a_66003_25280.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X627 a_28220_11501.t9 a_27762_11446.t28 a_27962_11501.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X628 vdd a_34044_31208.t96 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X629 a_64051_26022.t0 RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X630 a_65427_26048.t2 a_65077_26048.t2 a_65332_26048.t3 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X631 vdd a_34044_31208.t97 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X632 a_17685_3840.t9 vinit vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=1e+06u
X633 a_23145_17217.t4 Fvco.t31 a_22887_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X634 a_28994_17218.t5 a_26368_16652.t26 a_28736_17218.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X635 a_28220_11501.t8 a_27762_11446.t29 a_27962_11501.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X636 a_42782_16060.t6 vbiasot.t4 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=4e+06u
X637 vdd a_51138_19904.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X638 a_25815_17217.t12 a_23436_16644.t28 a_25557_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X639 a_23403_11500.t12 a_14266_8900.t36 a_23145_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X640 a_28220_17218.t10 a_26368_16652.t27 a_27962_17218.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X641 vdd a_1026_45630.t97 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X642 vdd a_1026_45630.t98 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X643 a_25815_17217.t11 a_23436_16644.t29 a_25557_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X644 vdd a_34044_31208.t98 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X645 vctrl.t1 CLK_BY_4_IPH_BAR.t2 a_34044_31208.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X646 a_65992_26048.t1 a_64911_26048.t5 a_65645_26290.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X647 a_52052_20224.t1 a_56334_19906.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X648 a_28994_17218.t4 a_26368_16652.t28 a_28736_17218.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X649 a_42550_16062.t2 Fvco_By4_QPH.t7 a_42574_15624.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X650 a_24177_5596.t9 a_14188_14050.t27 a_23919_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X651 vdd a_34044_31208.t99 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X652 vdd a_1026_45630.t99 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X653 a_23436_16644.t0 Fvco.t32 a_23178_16644.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X654 a_29510_17218.t3 a_26368_16652.t29 a_29252_17218.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X655 a_22629_5596.t4 a_14188_14050.t28 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X656 vdd a_34044_31208.t100 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X657 a_66003_25280.t3 a_65088_25280.t5 a_65656_25522.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X658 Vso6b.t0 a_14832_12082.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X659 a_28736_11501.t6 a_27762_11446.t30 a_28478_11501.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X660 gnd a_17685_3840.t42 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X661 vdd a_34044_31208.t101 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X662 a_4314_11660.t0 a_4226_11612.t3 a_4314_11564.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X663 a_29510_17218.t2 a_26368_16652.t30 a_29252_17218.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X664 gnd a_17685_3840.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X665 a_65343_25280.t1 CLK_BY_4_IPH_BAR gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X666 a_28736_11501.t5 a_27762_11446.t31 a_28478_11501.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X667 a_23919_5596.t1 a_14188_14050.t29 a_23661_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X668 vdd a_34044_31208.t102 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X669 vdd a_1026_45630.t100 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X670 vdd a_1026_45630.t101 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X671 a_28478_11501.t10 a_27762_11446.t32 a_28220_11501.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X672 a_24177_5596.t8 a_14188_14050.t30 a_23919_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X673 vdd a_1026_45630.t102 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X674 vdd a_1026_45630.t103 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X675 vdd a_1026_45630.t104 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X676 a_23414_5032.t1 a_14188_14050.t31 a_17685_3840.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X677 vdd vinit a_17685_3840.t8 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51683e+11p pd=1.09597e+06u as=0p ps=0u w=1e+06u l=1e+06u
X678 a_28736_17218.t12 a_26368_16652.t31 a_28478_17218.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X679 gnd a_17685_3840.t44 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X680 a_28736_5597.t6 a_26036_4988.t32 a_28478_5597.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X681 vdd a_1026_45630.t105 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X682 gnd a_17685_3840.t45 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X683 gnd a_17685_3840.t46 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X684 vdd a_34044_31208.t103 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X685 vdd a_1026_45630.t106 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X686 a_26331_11500.t3 a_25099_11445.t33 a_26073_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X687 vdd a_1026_45630.t107 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X688 vdd a_34044_31208.t104 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X689 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=7.58416e+11p pd=5.47985e+06u as=7.58416e+11p ps=5.47985e+06u w=5e+06u l=1e+06u
X690 a_23156_5032.t4 a_14188_14050.t32 a_24177_5596.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X691 vdd a_34044_31208.t105 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X692 vdd a_34044_31208.t106 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X693 vdd a_1026_45630.t108 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X694 vdd a_34044_31208.t107 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X695 a_28736_17218.t1 a_26368_16652.t32 a_28478_17218.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X696 a_27962_5597.t3 a_26036_4988.t33 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X697 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X698 vdd a_1026_45630.t109 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X699 vdd a_34044_31208.t108 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X700 vdd a_1026_45630.t110 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X701 a_4314_11756.t0 a_4288_11726.t3 a_4314_11660.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X702 a_23145_5596.t9 a_14188_14050.t33 a_22887_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X703 a_28478_5597.t13 a_26036_4988.t34 a_28220_5597.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X704 vdd a_34044_31208.t109 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X705 a_26331_11500.t2 a_25099_11445.t34 a_26073_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X706 a_23661_5596.t3 a_14188_14050.t34 a_23403_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X707 vdd a_1026_45630.t111 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X708 a_25778_4988.t5 a_23414_5032.t30 a_26847_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X709 vdd a_34044_31208.t110 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X710 a_28994_17218.t3 a_26368_16652.t33 a_28736_17218.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X711 a_26331_11500.t1 a_25099_11445.t35 a_26073_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X712 z.t4 a_51334_14126.t7 a_51276_14152.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X713 a_28578_5014.t3 a_26036_4988.t35 a_29510_5597.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X714 a_23145_17217.t3 Fvco.t33 a_22887_17217.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X715 a_23308_802.t1 Fvco.t34 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X716 vdd a_34044_31208.t111 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X717 a_28994_17218.t2 a_26368_16652.t34 a_28736_17218.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X718 a_26331_11500.t0 a_25099_11445.t36 a_26073_11500.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X719 a_23145_17217.t2 Fvco.t35 a_22887_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X720 a_42782_16060.t2 Fvco_By4_QPH_bar.t5 a_43010_16058.t0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X721 a_27962_5597.t2 a_26036_4988.t36 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X722 vdd a_34044_31208.t112 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X723 a_28220_17218.t9 a_26368_16652.t35 a_27962_17218.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X724 vdd a_34044_31208.t113 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X725 a_65343_25280.t2 CLK_BY_4_IPH_BAR vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X726 CLK_BY_4_IPH a_66178_25254.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X727 a_26331_17217.t3 a_23436_16644.t30 a_26073_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X728 a_23403_5596.t8 a_14188_14050.t35 a_23145_5596.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X729 vdd a_34044_31208.t114 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X730 vdd a_1026_45630.t112 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X731 a_23178_16644.t4 Fvco.t36 a_24177_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X732 a_28220_17218.t8 a_26368_16652.t36 a_27962_17218.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X733 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X734 a_22887_5596.t3 a_14188_14050.t36 a_22629_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X735 gnd a_17685_3840.t47 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X736 a_23661_5596.t2 a_14188_14050.t37 a_23403_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X737 vdd a_1026_45630.t113 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X738 a_26847_5596.t12 a_23414_5032.t31 a_26589_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X739 vdd Vso8b.t3 a_4226_11612.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X740 a_24177_5596.t7 a_14188_14050.t38 a_23919_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X741 vdd a_34044_31208.t115 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X742 a_65992_26048.t0 a_65077_26048.t3 a_65645_26290.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X743 a_28220_5597.t4 a_26036_4988.t37 a_27962_5597.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X744 vdd a_34044_31208.t116 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X745 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=7.58416e+11p pd=5.47985e+06u as=7.58416e+11p ps=5.47985e+06u w=5e+06u l=1e+06u
X746 a_65332_26048.t1 Fvco_By4_QPH.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X747 a_46856_19268.t1 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X748 a_23414_5032.t0 a_14188_14050.t31 a_23156_5032.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X749 a_22629_5596.t3 a_14188_14050.t39 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X750 a_26847_11500.t2 a_25099_11445.t37 a_26589_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X751 a_29510_5597.t8 a_26036_4988.t38 a_29252_5597.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X752 vdd Vso6b.t3 a_4288_11726.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X753 a_46856_21176.t0 a_51138_20858.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X754 a_26073_5596.t10 a_23414_5032.t32 a_25815_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X755 vdd a_34044_31208.t117 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X756 a_26847_11500.t1 a_25099_11445.t38 a_26589_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X757 a_28994_5597.t2 a_26036_4988.t39 a_28736_5597.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X758 vdd a_1026_45630.t114 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X759 a_26589_11500.t4 a_25099_11445.t39 a_26331_11500.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X760 a_51826_16054.t1 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X761 a_26036_4988.t0 a_23414_5032.t14 a_25778_4988.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X762 a_26589_5596.t1 a_23414_5032.t33 a_26331_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X763 a_28736_17218.t0 a_26368_16652.t37 a_28478_17218.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X764 gnd a_56334_20860.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X765 vdd a_1026_45630.t115 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X766 a_26847_17217.t5 a_23436_16644.t31 a_26589_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X767 a_28736_17218.t6 a_26368_16652.t38 a_28478_17218.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X768 a_14266_8900.t0 a_25099_11445.t15 a_17685_3840.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X769 a_23661_11500.t10 a_14266_8900.t37 a_23403_11500.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X770 a_25815_5596.t3 a_23414_5032.t34 a_25557_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X771 a_51636_13108.t0 Fvco_By4_QPH_bar.t6 a_51276_14152.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X772 a_28736_5597.t1 a_26036_4988.t40 a_28478_5597.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X773 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X774 a_29252_5597.t7 a_26036_4988.t41 a_28994_5597.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X775 vdd a_1026_45630.t116 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X776 vdd a_34044_31208.t118 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X777 bb.t4 Fvco_By4_QPH.t9 a_47760_15642.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X778 a_26073_5596.t9 a_23414_5032.t35 a_25815_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X779 vdd a_1026_45630.t117 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X780 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X781 vdd a_34044_31208.t119 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X782 a_38070_8852.t0 a_25099_11445.t40 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X783 vdd a_1026_45630.t118 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X784 vdd Vso2b.t3 a_4226_12188.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X785 a_23156_5032.t3 a_14188_14050.t40 a_24177_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X786 vdd a_34044_31208.t120 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X787 a_26110_16652.t3 a_23436_16644.t32 a_26847_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X788 vdd a_1026_45630.t119 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X789 a_23661_11500.t9 a_14266_8900.t38 a_23403_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X790 a_27962_5597.t1 a_26036_4988.t42 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X791 a_23661_11500.t8 a_14266_8900.t39 a_23403_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X792 vdd a_1026_45630.t120 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X793 vdd a_34044_31208.t121 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X794 a_28438_10874.t4 a_27762_11446.t33 a_29510_11501.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X795 a_55602_11692.t0 Fvco_By4_QPH_bar.t7 a_50320_14126.t0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X796 gnd a_17685_3840.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X797 a_28478_5597.t12 a_26036_4988.t43 a_28220_5597.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X798 a_25557_5596.t7 a_23414_5032.t36 a_25299_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X799 a_26331_5596.t7 a_23414_5032.t37 a_26073_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X800 a_23661_11500.t7 a_14266_8900.t40 a_23403_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X801 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X802 a_23661_5596.t1 a_14188_14050.t41 a_23403_5596.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X803 vdd a_34044_31208.t122 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X804 vdd Vso3b.t4 a_4226_11996.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X805 a_26073_17217.t0 a_23436_16644.t33 a_25815_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X806 a_27762_11446.t0 a_26368_16652.t24 a_28622_16652.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X807 gnd a_17685_3840.t49 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X808 a_25778_4988.t4 a_23414_5032.t38 a_26847_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X809 vdd a_1026_45630.t121 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X810 vdd a_34044_31208.t123 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X811 vdd a_1026_45630.t122 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X812 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X813 a_57726_5786.t2 a_57726_5786.t1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.06485e+11p ps=5.25039e+06u w=3e+06u l=1e+06u
X814 vdd a_65645_26290.t4 a_65535_26414.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X815 a_8752_10532.t0 Vso7b.t5 a_4226_11612.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X816 a_23661_17217.t10 Fvco.t37 a_23403_17217.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X817 vdd a_34044_31208.t124 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X818 aa.t3 Fvco_By4_QPH.t10 a_47968_16078.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X819 vdd a_34044_31208.t125 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X820 a_4314_12140.t0 a_4288_12110.t3 a_4314_12044.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X821 a_26331_17217.t2 a_23436_16644.t34 a_26073_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X822 a_28438_10874.t3 a_27762_11446.t34 a_29510_11501.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X823 a_56602_11692.t7 a_51636_13108.t10 a_52052_20860.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X824 a_25557_11500.t8 a_25099_11445.t41 a_25299_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X825 vdd a_34044_31208.t126 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X826 vdd a_34044_31208.t127 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X827 a_62961_26048.t1 a_62795_26048.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.70773e+10p ps=701421u w=640000u l=150000u
X828 gnd a_17685_3840.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X829 a_26331_17217.t1 a_23436_16644.t35 a_26073_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X830 a_28438_10874.t2 a_27762_11446.t35 a_29510_11501.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X831 vdd a_34044_31208.t128 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X832 vdd a_1026_45630.t123 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X833 vdd a_1026_45630.t124 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X834 a_25557_11500.t7 a_25099_11445.t42 a_25299_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X835 Fvco.t1 a_26036_4988.t20 a_17685_3840.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X836 a_25299_5596.t1 a_23414_5032.t39 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X837 vdd a_34044_31208.t129 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X838 vdd a_1026_45630.t125 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X839 a_23403_11500.t9 a_14266_8900.t41 a_23145_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X840 a_28438_10874.t1 a_27762_11446.t36 a_29510_11501.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X841 a_55602_11692.t1 Fvco_By4_QPH_bar.t8 a_51334_14126.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X842 a_25299_11500.t4 a_25099_11445.t43 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X843 vdd a_66178_25254.t4 a_66742_25280.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=9.70773e+10p pd=701421u as=0p ps=0u w=640000u l=150000u
X844 a_26847_5596.t11 a_23414_5032.t40 a_26589_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X845 vdd a_1026_45630.t126 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X846 vdd a_34044_31208.t130 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X847 a_28622_16652.t2 a_26368_16652.t39 a_29510_17218.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X848 a_25557_17217.t3 a_23436_16644.t36 a_25299_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X849 a_24177_11500.t2 a_14266_8900.t42 a_23919_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X850 a_28220_5597.t3 a_26036_4988.t44 a_27962_5597.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X851 vdd a_1026_45630.t127 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X852 vdd a_34044_31208.t131 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X853 a_26690_784.t0 a_23414_5032.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X854 vdd a_1026_45630.t128 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X855 vdd a_34044_31208.t132 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X856 a_29252_11501.t9 a_27762_11446.t37 a_28994_11501.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X857 a_24177_11500.t1 a_14266_8900.t43 a_23919_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X858 a_23403_11500.t8 a_14266_8900.t44 a_23145_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X859 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X860 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X861 vdd a_1026_45630.t129 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X862 a_29252_11501.t8 a_27762_11446.t38 a_28994_11501.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X863 a_55602_11692.t10 a_51041_13108.t10 a_52052_20860.t16 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X864 a_26073_5596.t8 a_23414_5032.t42 a_25815_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X865 a_23403_11500.t11 a_14266_8900.t45 a_23145_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X866 vdd a_1026_45630.t130 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X867 a_54966_3580.t1 a_49874_4150.t0 a_53308_3580.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.83e+06u l=8e+06u
X868 vdd a_1026_45630.t131 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X869 a_24177_17217.t6 Fvco.t38 a_23919_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X870 a_23403_11500.t10 a_14266_8900.t46 a_23145_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X871 a_25815_17217.t10 a_23436_16644.t37 a_25557_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X872 a_47760_15642.t0 Fvco_By4_QPH_bar.t9 bb.t0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X873 a_26589_5596.t4 a_23414_5032.t43 a_26331_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X874 vdd a_1026_45630.t132 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X875 vdd a_34044_31208.t133 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X876 a_63216_26048.t3 CLK_BY_2_BAR.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X877 a_26847_17217.t4 a_23436_16644.t38 a_26589_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X878 a_14188_14050.t1 a_14266_8900.t47 a_23160_10936.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X879 vdd a_34044_31208.t134 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X880 gnd a_4226_12188.t4 a_4314_12140.t1 gnd sky130_fd_pr__nfet_01v8 ad=7.63003e+11p pd=5.67042e+06u as=0p ps=0u w=3.24e+06u l=150000u
X881 vdd Vso5b.t4 a_4226_11804.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X882 a_29252_17218.t3 a_26368_16652.t40 a_28994_17218.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X883 a_23403_17217.t10 Fvco.t39 a_23145_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X884 a_26847_17217.t3 a_23436_16644.t39 a_26589_17217.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X885 a_28478_11501.t9 a_27762_11446.t39 a_28220_11501.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X886 a_51334_14126.t2 Fvco_By4_QPH.t11 a_55602_11692.t6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X887 vdd a_34044_31208.t135 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X888 a_62961_26048.t0 a_62795_26048.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X889 vdd a_64051_26022.t5 a_64615_26048.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=9.70773e+10p pd=701421u as=0p ps=0u w=640000u l=150000u
X890 gnd a_17685_3840.t51 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X891 vdd a_1026_45630.t133 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X892 vdd a_1026_45630.t134 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X893 vdd a_66178_25254.t5 a_66165_25646.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X894 Vso2b.t1 a_28790_25040.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X895 a_65700_25280.t1 a_65656_25522.t5 a_65534_25280.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X896 vdd a_34044_31208.t136 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X897 a_29252_17218.t2 a_26368_16652.t41 a_28994_17218.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X898 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X899 a_47760_15642.t1 Fvco_By4_QPH_bar.t10 aa.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X900 vdd a_34044_31208.t137 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X901 a_22972_23306.t1 a_23504_23306.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X902 a_28478_11501.t8 a_27762_11446.t40 a_28220_11501.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X903 a_50262_14152.t5 a_50320_14126.t6 a_50511_16072.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X904 vdd CLK_IN.t4 a_62795_26048.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=9.70773e+10p pd=701421u as=0p ps=0u w=640000u l=150000u
X905 CLK_BY_4_IPH_BAR a_66742_25280.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X906 a_23919_11500.t7 a_14266_8900.t48 a_23661_11500.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X907 a_28478_11501.t7 a_27762_11446.t41 a_28220_11501.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X908 vdd a_1026_45630.t135 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X909 a_65535_26414.t0 a_64911_26048.t6 a_65427_26048.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X910 vdd a_54468_7504.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X911 a_23919_11500.t10 a_14266_8900.t49 a_23661_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X912 a_28478_11501.t6 a_27762_11446.t42 a_28220_11501.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X913 a_26331_5596.t11 a_23414_5032.t44 a_26073_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X914 vdd a_1026_45630.t136 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X915 vdd a_1026_45630.t137 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X916 a_23661_17217.t9 Fvco.t40 a_23403_17217.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X917 vdd a_34044_31208.t138 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X918 a_22887_11500.t2 a_14266_8900.t50 a_22629_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X919 a_47968_16078.t0 Fvco_By4_QPH_bar.t11 bb.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X920 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X921 vdd a_1026_45630.t138 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X922 Vso1b.t0 a_24410_25128.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X923 a_28478_17218.t9 a_26368_16652.t42 a_28220_17218.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X924 a_23661_17217.t8 Fvco.t41 a_23403_17217.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X925 a_23919_17217.t13 Fvco.t42 a_23661_17217.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X926 a_22887_11500.t1 a_14266_8900.t51 a_22629_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X927 vdd a_1026_45630.t139 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X928 a_42550_16062.t3 Fvco_By4_QPH.t12 a_42782_16060.t5 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X929 vdd a_34044_31208.t139 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X930 vdd a_34044_31208.t140 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X931 a_22887_17217.t0 Fvco.t43 a_22629_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X932 a_52052_20860.t3 a_51636_13108.t11 a_56602_11692.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X933 Vso4b.t1 a_38070_8852.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X934 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X935 CLK_BY_2.t0 a_64051_26022.t6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X936 a_28622_16652.t1 a_26368_16652.t43 a_29510_17218.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X937 a_23145_5596.t8 a_14188_14050.t42 a_22887_5596.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X938 gnd RESET a_65700_25280.t0 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X939 gnd a_66178_25254.t6 a_66112_25280.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X940 a_25557_17217.t2 a_23436_16644.t40 a_25299_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X941 a_51532_4150.t0 a_49932_4124.t3 a_49874_4150.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.28e+06u l=8e+06u
X942 a_64725_25280.t1 CLK_BY_2_BAR.t7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X943 vdd a_4288_11534.t4 vout.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X944 a_28622_16652.t0 a_26368_16652.t44 a_29510_17218.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X945 vdd a_1026_45630.t140 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X946 CLK_BY_4_IPH.t0 a_66178_25254.t7 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X947 a_17685_3840.t16 vctrl.t4 a_22972_23306.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X948 a_25557_17217.t1 a_23436_16644.t41 a_25299_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X949 vdd a_34044_31208.t141 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X950 gnd CLK_IN.t5 a_62795_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X951 vdd a_34044_31208.t142 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X952 a_23145_17217.t1 Fvco.t44 a_22887_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X953 a_24177_17217.t5 Fvco.t45 a_23919_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X954 vdd a_1026_45630.t141 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X955 gnd a_17685_3840.t52 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X956 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=7.58416e+11p pd=5.47985e+06u as=7.58416e+11p ps=5.47985e+06u w=5e+06u l=1e+06u
X957 vdd a_34044_31208.t143 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X958 a_24177_17217.t4 Fvco.t46 a_23919_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X959 gnd a_17685_3840.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X960 vdd a_1026_45630.t142 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X961 a_29252_17218.t1 a_26368_16652.t45 a_28994_17218.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X962 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X963 vdd a_34044_31208.t144 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X964 a_65645_26290.t2 a_65427_26048.t5 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.27414e+11p ps=920615u w=840000u l=150000u
X965 a_23403_17217.t9 Fvco.t47 a_23145_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X966 a_52052_20860.t11 a_51041_13108.t11 a_55602_11692.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X967 a_22887_5596.t2 a_14188_14050.t43 a_22629_5596.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X968 vdd a_1026_45630.t143 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X969 vdd a_34044_31208.t145 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X970 a_29252_17218.t0 a_26368_16652.t46 a_28994_17218.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X971 vdd a_34044_31208.t146 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X972 vdd a_34044_31208.t147 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X973 a_23403_17217.t8 Fvco.t48 a_23145_17217.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X974 a_26589_11500.t1 a_25099_11445.t44 a_26331_11500.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X975 a_22629_11500.t1 a_14266_8900.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X976 a_24177_5596.t6 a_14188_14050.t44 a_23919_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X977 vdd a_1026_45630.t144 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X978 vdd a_34044_31208.t148 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X979 a_22629_11500.t0 a_14266_8900.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X980 vdd a_1026_45630.t145 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X981 a_50511_16072.t7 a_42550_16062.t5 a_47968_16078.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X982 vdd a_34044_31208.t149 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X983 vdd a_1026_45630.t146 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X984 vdd a_1026_45630.t147 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X985 vdd a_51138_20858.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X986 gnd a_17685_3840.t54 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X987 vdd a_1026_45630.t148 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X988 vdd a_1026_45630.t149 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X989 vdd a_34044_31208.t150 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X990 a_22629_17217.t2 Fvco.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X991 Fvco_By4_QPH.t1 a_66731_26048.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53072e+11p ps=1.13758e+06u w=650000u l=150000u
X992 Vso6b.t1 a_14832_12082.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X993 vdd Vso4b.t3 a_4226_11996.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X994 a_26589_11500.t0 a_25099_11445.t45 a_26331_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X995 a_50511_16072.t2 a_50320_14126.t7 a_50262_14152.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X996 a_56602_11692.t5 a_51636_13108.t12 a_52052_20860.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X997 a_51276_14152.t2 Fvco_By4_QPH.t13 a_51041_13108.t2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X998 a_28994_5597.t1 a_26036_4988.t45 a_28736_5597.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X999 a_26589_11500.t3 a_25099_11445.t46 a_26331_11500.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1000 vdd a_34044_31208.t151 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1001 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1002 vdd a_34044_31208.t152 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1003 vdd a_1026_45630.t150 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1004 vdd a_1026_45630.t151 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1005 a_26589_11500.t2 a_25099_11445.t47 a_26331_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1006 vdd a_1026_45630.t152 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1007 a_28478_17218.t8 a_26368_16652.t47 a_28220_17218.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1008 vdd a_34044_31208.t153 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1009 vdd a_1026_45630.t153 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1010 a_34044_31208.t3 CLK_BY_4_IPH.t4 vctrl.t2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1011 vdd Vso1b.t4 a_4226_12188.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1012 a_26589_17217.t5 a_23436_16644.t42 a_26331_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1013 a_23919_17217.t12 Fvco.t50 a_23661_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1014 a_28478_17218.t7 a_26368_16652.t48 a_28220_17218.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1015 a_28994_11501.t13 a_27762_11446.t43 a_28736_11501.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1016 vdd a_34044_31208.t154 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1017 a_56602_11692.t1 Fvco_By4_QPH_bar.t12 a_51334_14126.t1 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1018 a_63419_26414.t0 a_62795_26048.t5 a_63311_26048.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1019 a_23919_17217.t2 Fvco.t51 a_23661_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1020 a_43010_16058.t2 Fvco_By4_QPH.t14 a_42782_16060.t4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1021 vdd a_1026_45630.t154 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1022 vdd a_1026_45630.t155 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1023 a_55602_11692.t4 a_51041_13108.t12 a_52052_20860.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1024 vctrl.t0 CLK_BY_4_IPH_BAR.t3 a_1026_45630.t0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1025 a_24410_25128.t0 a_23436_16644.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X1026 a_63876_26048.t1 a_62795_26048.t6 a_63529_26290.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1027 a_22887_17217.t5 Fvco.t52 a_22629_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1028 a_53292_4814.t0 a_49874_4150.t0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.01433e+11p ps=2.24017e+06u w=1.28e+06u l=8e+06u
X1029 a_27962_5597.t0 a_26036_4988.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1030 gnd a_66167_26022.t7 a_66101_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X1031 gnd RESET a_65689_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X1032 a_22887_17217.t12 Fvco.t53 a_22629_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1033 vdd a_1026_45630.t156 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1034 gnd a_17685_3840.t55 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1035 a_22629_5596.t2 a_14188_14050.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1036 gnd a_17685_3840.t56 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1037 a_23145_5596.t13 a_14188_14050.t46 a_22887_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1038 vdd a_34044_31208.t155 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1039 vdd a_34044_31208.t156 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1040 a_63529_26290.t3 a_63311_26048.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.50717e+11p ps=1.12008e+06u w=640000u l=150000u
X1041 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.35495e+11p pd=1.75013e+06u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1042 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.29693e+12p pd=2.45018e+07u as=3.29693e+12p ps=2.45018e+07u w=1.4e+07u l=1e+06u
X1043 a_23661_5596.t0 a_14188_14050.t47 a_23403_5596.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1044 vdd a_1026_45630.t157 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1045 a_28790_25040.t0 a_26368_16652.t49 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X1046 a_25299_11500.t3 a_25099_11445.t48 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1047 vdd a_1026_45630.t158 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1048 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1049 Vso8b.t0 a_30384_802.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=9.89078e+10p ps=735055u w=420000u l=150000u
X1050 vdd Vso2b.t4 a_4288_12110.t0 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1051 a_46856_19268.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1052 vdd a_34044_31208.t157 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1053 vdd Vso4b.t4 a_4288_11918.t1 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1054 a_56602_11692.t4 a_51636_13108.t13 a_52052_20860.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1055 gnd a_17685_3840.t57 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1056 a_42782_16060.t1 bb.t5 a_44752_16348.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1057 vdd a_34044_31208.t158 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1058 a_64051_26022.t1 a_63876_26048.t5 a_64230_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1059 a_8748_11114.t0 Vso6b.t4 a_4288_11726.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1060 a_26331_17217.t0 a_23436_16644.t44 a_26073_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1061 a_22629_5596.t1 a_14188_14050.t48 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1062 a_28736_5597.t0 a_26036_4988.t47 a_28478_5597.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1063 vdd a_34044_31208.t159 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1064 a_25299_11500.t2 a_25099_11445.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1065 a_22887_5596.t1 a_14188_14050.t49 a_22629_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1066 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1067 vdd a_1026_45630.t159 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1068 a_25299_11500.t1 a_25099_11445.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1069 a_23919_5596.t0 a_14188_14050.t50 a_23661_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1070 vdd a_34044_31208.t160 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1071 a_28736_11501.t4 a_27762_11446.t44 a_28478_11501.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1072 vbiasot.t0 a_51532_4150.t6 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=8.1909e+10p ps=591824u w=540000u l=8e+06u
X1073 a_27962_11501.t1 a_27762_11446.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1074 a_25299_11500.t0 a_25099_11445.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1075 vbiasbuffer.t1 vbiasbuffer.t0 a_54468_7504.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1076 a_23156_5032.t2 a_14188_14050.t51 a_24177_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1077 vdd a_34044_31208.t161 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1078 a_14188_14050.t0 a_14266_8900.t47 a_17685_3840.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1079 a_27962_11501.t0 a_27762_11446.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1080 a_55602_11692.t2 a_51041_13108.t13 a_52052_20860.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=1e+06u
X1081 a_51334_14126.t3 Fvco_By4_QPH.t15 a_56602_11692.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1082 vdd a_34044_31208.t162 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1083 a_25299_17217.t2 a_23436_16644.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1084 a_22629_17217.t1 Fvco.t54 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1085 gnd a_17685_3840.t58 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1086 vdd a_1026_45630.t160 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1087 a_42574_15624.t5 aa.t5 a_44752_16348.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1088 vdd a_1026_45630.t161 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1089 a_28736_5597.t5 a_26036_4988.t48 a_28478_5597.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1090 a_26073_5596.t7 a_23414_5032.t45 a_25815_5596.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1091 a_24410_25128.t1 a_23436_16644.t12 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X1092 vdd a_4288_11726.t4 vout.t9 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1093 a_14832_12082.t0 a_14188_14050.t52 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X1094 a_22629_17217.t0 Fvco.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1095 a_50128_8156.t0 a_54410_8156.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1096 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1097 a_28994_5597.t0 a_26036_4988.t49 a_28736_5597.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1098 a_28478_5597.t10 a_26036_4988.t50 a_28220_5597.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1099 vdd a_34044_31208.t163 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1100 a_23160_10936.t2 a_14266_8900.t54 a_24177_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1101 a_42574_15624.t1 Fvco_By4_QPH_bar.t13 a_43010_16058.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1102 a_17685_3840.t7 vinit vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=1e+06u
X1103 a_27962_17218.t3 a_26368_16652.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1104 a_54966_2992.t0 a_49874_4150.t0 a_53308_2992.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.35e+06u l=8e+06u
X1105 a_25778_4988.t3 a_23414_5032.t46 a_26847_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1106 a_25099_11445.t0 a_27762_11446.t11 a_17685_3840.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1107 a_23160_10936.t1 a_14266_8900.t55 a_24177_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1108 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1109 vdd a_1026_45630.t162 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1110 a_22972_23306.t3 vctrl.t5 a_17685_3840.t15 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1111 a_23156_5032.t1 a_14188_14050.t53 a_24177_5596.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1112 vdd a_34044_31208.t164 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1113 vdd a_1026_45630.t163 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1114 vdd a_34044_31208.t165 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1115 vdd a_34044_31208.t166 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1116 vdd a_1026_45630.t164 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1117 a_17685_3840.t14 vctrl.t6 a_22972_23306.t2 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1118 a_26589_17217.t4 a_23436_16644.t46 a_26331_17217.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1119 vdd a_1026_45630.t165 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1120 a_8740_12844.t1 Vso3b.t5 a_4226_11996.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1121 a_4314_11468.t1 a_4226_11420.t4 vout.t5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X1122 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1123 a_66154_26414.t1 a_65077_26048.t4 a_65992_26048.t2 vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1124 a_27762_11446.t1 a_26368_16652.t24 a_17685_3840.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1125 a_26589_17217.t13 a_23436_16644.t47 a_26331_17217.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1126 a_38070_8852.t1 a_25099_11445.t52 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.34258e+10p ps=602784u w=550000u l=8e+06u
X1127 a_23178_16644.t3 Fvco.t56 a_24177_17217.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1128 a_27962_17218.t2 a_26368_16652.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1129 a_28478_5597.t9 a_26036_4988.t51 a_28220_5597.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1130 vdd a_1026_45630.t166 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1131 vdd a_34044_31208.t167 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1132 a_22972_23306.t0 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X1133 a_51041_13108.t1 Fvco_By4_QPH_bar.t14 a_50262_14152.t0 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1134 a_25778_4988.t2 a_23414_5032.t47 a_26847_5596.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1135 vdd a_34044_31208.t168 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1136 a_26847_5596.t10 a_23414_5032.t48 a_26589_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1137 vdd a_1026_45630.t167 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1138 a_32948_24994.t0 a_27762_11446.t47 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=150000u
X1139 a_28578_5014.t2 a_26036_4988.t52 a_29510_5597.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1140 vdd a_34044_31208.t169 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1141 vdd a_1026_45630.t168 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1142 vdd a_1026_45630.t169 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1143 a_63419_26414.t1 RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X1144 a_28220_5597.t2 a_26036_4988.t53 a_27962_5597.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1145 vdd a_1026_45630.t170 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1146 vdd a_1026_45630.t171 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1147 a_22629_5596.t0 a_14188_14050.t54 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1148 a_55602_11692.t13 vbiasob.t4 a_51138_21494.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X1149 a_23403_5596.t7 a_14188_14050.t55 a_23145_5596.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1150 vdd a_1026_45630.t172 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1151 vdd a_34044_31208.t170 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1152 vdd a_34044_31208.t171 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1153 vdd a_34044_31208.t172 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1154 vdd a_1026_45630.t173 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1155 vdd a_34044_31208.t173 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1156 vdd a_1026_45630.t174 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1157 vdd a_4226_11612.t4 vout.t8 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1158 a_23661_17217.t7 Fvco.t57 a_23403_17217.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1159 a_51041_13108.t0 Fvco_By4_QPH_bar.t15 a_51276_14152.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1160 a_26847_5596.t6 a_23414_5032.t49 a_26589_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1161 vdd a_34044_31208.t174 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1162 a_26589_5596.t3 a_23414_5032.t50 a_26331_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1163 a_28220_5597.t1 a_26036_4988.t54 a_27962_5597.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1164 vdd a_1026_45630.t175 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1165 vdd a_1026_45630.t176 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1166 vdd a_64051_26022.t7 a_64038_26414.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X1167 a_4314_11852.t1 a_4226_11804.t3 a_4314_11756.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X1168 a_26016_10878.t1 a_25099_11445.t53 a_26847_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1169 vdd a_1026_45630.t177 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1170 gnd a_66178_25254.t8 a_66742_25280.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X1171 a_26016_10878.t0 a_25099_11445.t54 a_26847_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1172 a_28736_5597.t4 a_26036_4988.t55 a_28478_5597.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1173 a_29510_5597.t7 a_26036_4988.t56 a_29252_5597.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1174 aa.t2 vbiasbuffer.t4 a_50032_16080.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1175 a_26847_11500.t0 a_25099_11445.t55 a_26589_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1176 a_51636_13108.t1 Fvco_By4_QPH_bar.t16 a_50262_14152.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1177 vdd a_66003_25280.t4 a_66178_25254.t1 vdd sky130_fd_pr__pfet_01v8_hvt ad=6.3707e+10p pd=460307u as=0p ps=0u w=420000u l=150000u
X1178 a_8748_11692.t1 Vso5b.t5 a_4226_11804.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1179 a_26073_11500.t10 a_25099_11445.t56 a_25815_11500.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1180 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=7.58416e+11p pd=5.47985e+06u as=7.58416e+11p ps=5.47985e+06u w=5e+06u l=1e+06u
X1181 a_50262_14152.t3 Fvco_By4_QPH.t16 a_51636_13108.t3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1182 a_23156_5032.t0 a_14188_14050.t56 a_24177_5596.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1183 CLK_BY_2_BAR.t1 a_64615_26048.t3 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.51683e+11p ps=1.09597e+06u w=1e+06u l=150000u
X1184 a_8744_9386.t1 CLK_IN.t6 a_4226_11420.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1185 gnd a_17685_3840.t59 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1186 a_26589_5596.t6 a_23414_5032.t51 a_26331_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1187 vdd a_34044_31208.t175 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1188 a_26110_16652.t2 a_23436_16644.t48 a_26847_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1189 a_25299_17217.t1 a_23436_16644.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1190 a_26073_11500.t11 a_25099_11445.t57 a_25815_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1191 vdd a_34044_31208.t176 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1192 vdd a_1026_45630.t178 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1193 a_65427_26048.t0 a_64911_26048.t7 a_65332_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1194 vdd a_64725_25280.t5 a_64922_25280.t0 vdd sky130_fd_pr__pfet_01v8_hvt ad=9.70773e+10p pd=701421u as=0p ps=0u w=640000u l=150000u
X1195 a_25299_17217.t0 a_23436_16644.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1196 gnd a_17685_3840.t60 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1197 vdd a_34044_31208.t177 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1198 a_44752_16348.t1 bb.t6 a_42782_16060.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1199 a_25815_5596.t2 a_23414_5032.t52 a_25557_5596.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1200 a_27962_17218.t1 a_26368_16652.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1201 gnd a_17685_3840.t61 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1202 a_28478_5597.t11 a_26036_4988.t57 a_28220_5597.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1203 a_26331_5596.t10 a_23414_5032.t53 a_26073_5596.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1204 vdd a_34044_31208.t178 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1205 a_66178_25254.t0 a_66003_25280.t5 a_66357_25280.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1206 gnd Vso8b.t4 a_8752_10532.t1 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X1207 a_29252_5597.t6 a_26036_4988.t58 a_28994_5597.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1208 a_26073_17217.t2 a_23436_16644.t51 a_25815_17217.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1209 a_27962_17218.t0 a_26368_16652.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1210 a_25778_4988.t1 a_23414_5032.t54 a_26847_5596.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1211 vdd a_1026_45630.t179 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1212 vdd a_34044_31208.t179 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1213 a_47760_15642.t5 a_43010_16058.t4 z.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1214 vdd a_34044_31208.t180 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1215 a_63529_26290.t1 a_63311_26048.t5 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=1.27414e+11p ps=920615u w=840000u l=150000u
X1216 vdd a_1026_45630.t180 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1217 a_23403_17217.t7 Fvco.t58 a_23145_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1218 vdd a_34044_31208.t181 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1219 vdd a_34044_31208.t182 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1220 a_4314_11948.t1 a_4288_11918.t4 a_4314_11852.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.24e+06u l=150000u
X1221 gnd a_17685_3840.t62 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1222 a_23178_16644.t2 Fvco.t59 a_24177_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1223 a_51532_4150.t3 a_49874_4150.t0 a_54966_3580.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.83e+06u l=8e+06u
X1224 gnd CLK_BY_2_BAR.t8 a_64725_25280.t0 gnd sky130_fd_pr__nfet_01v8 ad=1.53072e+11p pd=1.13758e+06u as=0p ps=0u w=650000u l=150000u
X1225 vdd a_1026_45630.t181 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1226 a_23178_16644.t1 Fvco.t60 a_24177_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1227 a_25557_5596.t13 a_23414_5032.t55 a_25299_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1228 vdd a_1026_45630.t182 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1229 a_44752_16348.t0 aa.t6 a_42574_15624.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1230 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1231 a_26331_5596.t13 a_23414_5032.t56 a_26073_5596.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1232 vdd a_1026_45630.t183 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1233 gnd Vso6b.t5 a_8748_11692.t0 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X1234 a_28994_11501.t1 a_27762_11446.t48 a_28736_11501.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1235 a_26847_5596.t5 a_23414_5032.t57 a_26589_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1236 a_65332_26048.t2 Fvco_By4_QPH.t17 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X1237 a_25815_11500.t8 a_25099_11445.t58 a_25557_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1238 a_28220_5597.t0 a_26036_4988.t59 a_27962_5597.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1239 vdd a_1026_45630.t184 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1240 a_25815_11500.t7 a_25099_11445.t59 a_25557_11500.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1241 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1242 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1243 vdd a_1026_45630.t185 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1244 a_8748_9956.t1 Vso8b.t5 a_4288_11534.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1245 gnd a_17685_3840.t63 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1246 a_25557_11500.t6 a_25099_11445.t60 a_25299_11500.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1247 vdd a_34044_31208.t183 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1248 a_28994_11501.t0 a_27762_11446.t49 a_28736_11501.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1249 a_25299_5596.t0 a_23414_5032.t58 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=2.35495e+11p ps=1.75013e+06u w=1e+06u l=1e+06u
X1250 vdd a_34044_31208.t184 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1251 vdd a_34044_31208.t185 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1252 a_66178_25254.t2 RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X1253 a_28994_11501.t10 a_27762_11446.t50 a_28736_11501.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1254 vdd a_4288_12110.t4 vout.t2 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1255 a_25815_17217.t9 a_23436_16644.t52 a_25557_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1256 a_26589_5596.t5 a_23414_5032.t59 a_26331_5596.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1257 a_28994_11501.t11 a_27762_11446.t51 a_28736_11501.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1258 Vso8b.t1 a_30384_802.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.54828e+11p ps=1.84123e+06u w=1.68e+06u l=150000u
X1259 gnd a_66167_26022.t8 a_66731_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X1260 a_29510_11501.t8 a_27762_11446.t52 a_29252_11501.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1261 vdd a_34044_31208.t186 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1262 vdd a_34044_31208.t187 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1263 a_24177_11500.t0 a_14266_8900.t56 a_23919_11500.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1264 z.t0 a_43010_16058.t5 a_47760_15642.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1265 vdd a_34044_31208.t188 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1266 vdd a_1026_45630.t186 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1267 vdd a_1026_45630.t187 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1268 a_29510_11501.t7 a_27762_11446.t53 a_29252_11501.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1269 vdd a_34044_31208.t189 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1270 a_28994_17218.t1 a_26368_16652.t54 a_28736_17218.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1271 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1272 gnd a_17685_3840.t64 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.64846e+12p pd=1.22509e+07u as=1.64846e+12p ps=1.22509e+07u w=7e+06u l=8e+06u
X1273 a_29252_11501.t7 a_27762_11446.t54 a_28994_11501.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1274 a_42782_16060.t3 Fvco_By4_QPH_bar.t17 a_42550_16062.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1275 vdd a_34044_31208.t190 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1276 gnd a_64051_26022.t8 a_63985_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=9.89078e+10p pd=735055u as=0p ps=0u w=420000u l=150000u
X1277 vdd a_1026_45630.t188 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1278 vdd a_1026_45630.t189 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1279 a_26110_16652.t1 a_23436_16644.t53 a_26847_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1280 a_50320_14126.t3 Fvco_By4_QPH.t18 a_56602_11692.t2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1281 a_29510_17218.t1 a_26368_16652.t55 a_29252_17218.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1282 a_63985_26048.t0 a_62795_26048.t7 a_63876_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1283 a_26110_16652.t0 a_23436_16644.t54 a_26847_17217.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1284 vdd a_34044_31208.t191 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1285 vdd a_34044_31208.t192 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1286 vdd a_34044_31208.t193 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1287 a_28736_11501.t3 a_27762_11446.t55 a_28478_11501.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1288 a_50262_14152.t8 a_50320_14126.t8 a_50511_16072.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1289 vdd a_1026_45630.t190 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1290 vdd a_34044_31208.t194 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1291 a_66167_26022.t1 a_65992_26048.t5 a_66346_26048.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1292 vdd a_34044_31208.t195 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1293 vdd a_34044_31208.t196 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1294 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1295 a_26073_17217.t5 a_23436_16644.t55 a_25815_17217.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1296 a_51276_14152.t5 a_51334_14126.t8 z.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1297 vdd a_34044_31208.t197 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1298 vdd a_1026_45630.t191 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1299 a_26331_5596.t12 a_23414_5032.t60 a_26073_5596.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1300 a_26073_17217.t3 a_23436_16644.t56 a_25815_17217.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1301 vdd a_4226_11804.t4 vout.t7 vdd sky130_fd_pr__pfet_01v8 ad=2.54828e+11p pd=1.84123e+06u as=0p ps=0u w=1.68e+06u l=150000u
X1302 a_29510_17218.t0 a_26368_16652.t56 a_29252_17218.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1303 vdd a_1026_45630.t192 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1304 a_28736_11501.t2 a_27762_11446.t56 a_28478_11501.t2 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1305 vdd a_1026_45630.t193 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1306 a_65088_25280.t0 a_64922_25280.t7 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=9.70773e+10p ps=701421u w=640000u l=150000u
X1307 vdd a_34044_31208.t198 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1308 a_28736_11501.t1 a_27762_11446.t57 a_28478_11501.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1309 a_50511_16072.t0 a_50320_14126.t9 a_50262_14152.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1310 a_23919_5596.t2 a_14188_14050.t57 a_23661_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1311 vdd a_1026_45630.t194 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1312 a_28736_11501.t0 a_27762_11446.t58 a_28478_11501.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1313 vdd a_34044_31208.t199 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1314 a_23919_11500.t9 a_14266_8900.t57 a_23661_11500.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1315 vdd a_1026_45630.t195 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1316 vdd a_1026_45630.t196 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1317 a_8736_14034.t0 Vso1b.t5 a_4226_12188.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1318 vdd a_1026_45630.t197 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1319 a_65689_26048.t0 a_65645_26290.t5 a_65523_26048.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1320 a_28736_17218.t5 a_26368_16652.t57 a_28478_17218.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1321 a_23145_11500.t8 a_14266_8900.t58 a_22887_11500.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1322 a_23145_5596.t12 a_14188_14050.t58 a_22887_5596.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1323 a_63876_26048.t3 a_62961_26048.t5 a_63529_26290.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1324 a_23145_11500.t7 a_14266_8900.t59 a_22887_11500.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1325 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1326 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1327 a_65523_26048.t1 a_65077_26048.t5 a_65427_26048.t3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1328 gnd CLK_IN.t7 a_8748_9956.t0 gnd sky130_fd_pr__nfet_01v8 ad=1.74266e+11p pd=1.2951e+06u as=0p ps=0u w=740000u l=150000u
X1329 a_28220_11501.t7 a_27762_11446.t59 a_27962_11501.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1330 a_22887_11500.t0 a_14266_8900.t60 a_22629_11500.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1331 vdd a_1026_45630.t198 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1332 vdd a_1026_45630.t199 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1333 a_28220_11501.t6 a_27762_11446.t60 a_27962_11501.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1334 vdd a_1026_45630.t200 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1335 vdd a_34044_31208.t200 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1336 vdd a_1026_45630.t201 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1337 vdd a_34044_31208.t201 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1338 a_23145_17217.t0 Fvco.t61 a_22887_17217.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1339 a_63216_26048.t2 CLK_BY_2_BAR.t9 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=6.3707e+10p ps=460307u w=420000u l=150000u
X1340 vdd a_1026_45630.t202 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1341 a_25815_17217.t8 a_23436_16644.t57 a_25557_17217.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1342 z.t2 a_51334_14126.t9 a_51276_14152.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X1343 a_28220_17218.t7 a_26368_16652.t58 a_27962_17218.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1344 a_26589_17217.t12 a_23436_16644.t58 a_26331_17217.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1345 vdd a_34044_31208.t202 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1346 a_26368_16652.t0 a_23436_16644.t12 a_17685_3840.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1347 a_25815_17217.t7 a_23436_16644.t59 a_25557_17217.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1348 a_23145_5596.t0 a_14188_14050.t59 a_22887_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1349 vdd a_34044_31208.t203 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
X1350 a_8744_13422.t0 Vso2b.t5 a_4288_12110.t1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1351 aa.t4 Fvco_By4_QPH.t19 a_47760_15642.t3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X1352 a_22887_5596.t0 a_14188_14050.t60 a_22629_5596.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1353 a_8748_12270.t0 Vso4b.t5 a_4288_11918.t0 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1354 a_28994_17218.t0 a_26368_16652.t59 a_28736_17218.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1355 a_28578_5014.t1 a_26036_4988.t60 a_29510_5597.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1356 vdd a_1026_45630.t203 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.06178e+12p pd=7.67179e+06u as=1.06178e+12p ps=7.67179e+06u w=7e+06u l=8e+06u
C0 vdd Vso5b 5.20fF
C1 vdd CLK_IN 2.08fF
C2 vdd Vso3b 3.96fF
C3 vdd vbiasob 2.62fF
C4 vdd Vso4b 3.85fF
C5 CLK_IN Vso4b 26.23fF
C6 vdd Fvco_By4_QPH_bar 2.21fF
C7 Fvco_By4_QPH Fvco_By4_QPH_bar 16.00fF
C8 CLK_BY_4_IPH_BAR CLK_BY_4_IPH 11.02fF
C9 vdd vout 7.94fF
C10 vdd Vso7b 2.92fF
C11 vdd Vso6b 3.09fF
C12 vdd Fvco 4.89fF
C13 RESET Fvco_By4_QPH 2.21fF
C14 vdd CLK_BY_4_IPH_BAR 14.46fF
C15 Fvco_By4_QPH_bar bb 2.30fF
C16 Vso7b Vso8b 12.19fF
C17 vdd Vso2b 3.24fF
C18 aa bb 2.62fF
R0 a_34044_31208.n0 a_34044_31208.t3 16.252
R1 a_34044_31208.t1 a_34044_31208.n0 16.252
R2 a_34044_31208.n0 a_34044_31208.n204 1.906
R3 a_34044_31208.n204 a_34044_31208.n2 38.8
R4 a_34044_31208.n2 a_34044_31208.n13 0.514
R5 a_34044_31208.n2 a_34044_31208.n3 6.785
R6 a_34044_31208.n8 a_34044_31208.n14 1.97
R7 a_34044_31208.n14 a_34044_31208.n9 17.089
R8 a_34044_31208.n9 a_34044_31208.n10 7.911
R9 a_34044_31208.n13 a_34044_31208.n194 56.763
R10 a_34044_31208.n194 a_34044_31208.n203 7.74
R11 a_34044_31208.n203 a_34044_31208.t73 7.285
R12 a_34044_31208.n203 a_34044_31208.n202 14.37
R13 a_34044_31208.n202 a_34044_31208.t139 7.285
R14 a_34044_31208.n202 a_34044_31208.n201 14.37
R15 a_34044_31208.n201 a_34044_31208.t183 7.285
R16 a_34044_31208.n201 a_34044_31208.n200 14.37
R17 a_34044_31208.n200 a_34044_31208.t56 7.285
R18 a_34044_31208.n200 a_34044_31208.n199 14.395
R19 a_34044_31208.n199 a_34044_31208.t104 7.285
R20 a_34044_31208.n199 a_34044_31208.n198 14.37
R21 a_34044_31208.n198 a_34044_31208.t60 7.285
R22 a_34044_31208.n198 a_34044_31208.n197 14.37
R23 a_34044_31208.n197 a_34044_31208.t126 7.285
R24 a_34044_31208.n197 a_34044_31208.n196 14.37
R25 a_34044_31208.n196 a_34044_31208.t170 7.285
R26 a_34044_31208.n196 a_34044_31208.n195 15.728
R27 a_34044_31208.n195 a_34044_31208.t85 7.285
R28 a_34044_31208.n195 a_34044_31208.t151 21.655
R29 a_34044_31208.n194 a_34044_31208.n184 64.823
R30 a_34044_31208.n184 a_34044_31208.n193 7.74
R31 a_34044_31208.n193 a_34044_31208.t34 7.285
R32 a_34044_31208.n193 a_34044_31208.n192 14.37
R33 a_34044_31208.n192 a_34044_31208.t100 7.285
R34 a_34044_31208.n192 a_34044_31208.n191 14.37
R35 a_34044_31208.n191 a_34044_31208.t145 7.285
R36 a_34044_31208.n191 a_34044_31208.n190 14.37
R37 a_34044_31208.n190 a_34044_31208.t16 7.285
R38 a_34044_31208.n190 a_34044_31208.n189 14.395
R39 a_34044_31208.n189 a_34044_31208.t68 7.285
R40 a_34044_31208.n189 a_34044_31208.n188 14.37
R41 a_34044_31208.n188 a_34044_31208.t21 7.285
R42 a_34044_31208.n188 a_34044_31208.n187 14.37
R43 a_34044_31208.n187 a_34044_31208.t87 7.285
R44 a_34044_31208.n187 a_34044_31208.n186 14.37
R45 a_34044_31208.n186 a_34044_31208.t133 7.285
R46 a_34044_31208.n186 a_34044_31208.n185 15.728
R47 a_34044_31208.n185 a_34044_31208.t45 7.285
R48 a_34044_31208.n185 a_34044_31208.t113 21.655
R49 a_34044_31208.n184 a_34044_31208.n174 62.638
R50 a_34044_31208.n174 a_34044_31208.n183 7.74
R51 a_34044_31208.n183 a_34044_31208.t125 7.285
R52 a_34044_31208.n183 a_34044_31208.n182 14.37
R53 a_34044_31208.n182 a_34044_31208.t193 7.285
R54 a_34044_31208.n182 a_34044_31208.n181 14.37
R55 a_34044_31208.n181 a_34044_31208.t40 7.285
R56 a_34044_31208.n181 a_34044_31208.n180 14.37
R57 a_34044_31208.n180 a_34044_31208.t106 7.285
R58 a_34044_31208.n180 a_34044_31208.n179 14.395
R59 a_34044_31208.n179 a_34044_31208.t156 7.285
R60 a_34044_31208.n179 a_34044_31208.n178 14.37
R61 a_34044_31208.n178 a_34044_31208.t111 7.285
R62 a_34044_31208.n178 a_34044_31208.n177 14.37
R63 a_34044_31208.n177 a_34044_31208.t175 7.285
R64 a_34044_31208.n177 a_34044_31208.n176 14.37
R65 a_34044_31208.n176 a_34044_31208.t26 7.285
R66 a_34044_31208.n176 a_34044_31208.n175 15.728
R67 a_34044_31208.n175 a_34044_31208.t137 7.285
R68 a_34044_31208.n175 a_34044_31208.t203 21.655
R69 a_34044_31208.n174 a_34044_31208.n164 58.45
R70 a_34044_31208.n164 a_34044_31208.n173 7.74
R71 a_34044_31208.n173 a_34044_31208.t194 7.285
R72 a_34044_31208.n173 a_34044_31208.n172 14.37
R73 a_34044_31208.n172 a_34044_31208.t63 7.285
R74 a_34044_31208.n172 a_34044_31208.n171 14.37
R75 a_34044_31208.n171 a_34044_31208.t107 7.285
R76 a_34044_31208.n171 a_34044_31208.n170 14.37
R77 a_34044_31208.n170 a_34044_31208.t174 7.285
R78 a_34044_31208.n170 a_34044_31208.n169 14.395
R79 a_34044_31208.n169 a_34044_31208.t28 7.285
R80 a_34044_31208.n169 a_34044_31208.n168 14.37
R81 a_34044_31208.n168 a_34044_31208.t176 7.285
R82 a_34044_31208.n168 a_34044_31208.n167 14.37
R83 a_34044_31208.n167 a_34044_31208.t48 7.285
R84 a_34044_31208.n167 a_34044_31208.n166 14.37
R85 a_34044_31208.n166 a_34044_31208.t92 7.285
R86 a_34044_31208.n166 a_34044_31208.n165 15.728
R87 a_34044_31208.n165 a_34044_31208.t55 7.285
R88 a_34044_31208.n165 a_34044_31208.t120 21.655
R89 a_34044_31208.n164 a_34044_31208.n154 58.268
R90 a_34044_31208.n154 a_34044_31208.n163 7.74
R91 a_34044_31208.n163 a_34044_31208.t136 7.285
R92 a_34044_31208.n163 a_34044_31208.n162 14.37
R93 a_34044_31208.n162 a_34044_31208.t202 7.285
R94 a_34044_31208.n162 a_34044_31208.n161 14.37
R95 a_34044_31208.n161 a_34044_31208.t52 7.285
R96 a_34044_31208.n161 a_34044_31208.n160 14.37
R97 a_34044_31208.n160 a_34044_31208.t117 7.285
R98 a_34044_31208.n160 a_34044_31208.n159 14.395
R99 a_34044_31208.n159 a_34044_31208.t166 7.285
R100 a_34044_31208.n159 a_34044_31208.n158 14.37
R101 a_34044_31208.n158 a_34044_31208.t119 7.285
R102 a_34044_31208.n158 a_34044_31208.n157 14.37
R103 a_34044_31208.n157 a_34044_31208.t184 7.285
R104 a_34044_31208.n157 a_34044_31208.n156 14.37
R105 a_34044_31208.n156 a_34044_31208.t35 7.285
R106 a_34044_31208.n156 a_34044_31208.n155 15.728
R107 a_34044_31208.n155 a_34044_31208.t143 7.285
R108 a_34044_31208.n155 a_34044_31208.t14 21.655
R109 a_34044_31208.n154 a_34044_31208.n144 63.367
R110 a_34044_31208.n144 a_34044_31208.n153 7.74
R111 a_34044_31208.n153 a_34044_31208.t95 7.285
R112 a_34044_31208.n153 a_34044_31208.n152 14.37
R113 a_34044_31208.n152 a_34044_31208.t160 7.285
R114 a_34044_31208.n152 a_34044_31208.n151 14.37
R115 a_34044_31208.n151 a_34044_31208.t7 7.285
R116 a_34044_31208.n151 a_34044_31208.n150 14.37
R117 a_34044_31208.n150 a_34044_31208.t75 7.285
R118 a_34044_31208.n150 a_34044_31208.n149 14.395
R119 a_34044_31208.n149 a_34044_31208.t129 7.285
R120 a_34044_31208.n149 a_34044_31208.n148 14.37
R121 a_34044_31208.n148 a_34044_31208.t80 7.285
R122 a_34044_31208.n148 a_34044_31208.n147 14.37
R123 a_34044_31208.n147 a_34044_31208.t146 7.285
R124 a_34044_31208.n147 a_34044_31208.n146 14.37
R125 a_34044_31208.n146 a_34044_31208.t195 7.285
R126 a_34044_31208.n146 a_34044_31208.n145 15.728
R127 a_34044_31208.n145 a_34044_31208.t103 7.285
R128 a_34044_31208.n145 a_34044_31208.t173 21.655
R129 a_34044_31208.n144 a_34044_31208.n134 62.456
R130 a_34044_31208.n134 a_34044_31208.n143 7.74
R131 a_34044_31208.n143 a_34044_31208.t9 7.285
R132 a_34044_31208.n143 a_34044_31208.n142 14.37
R133 a_34044_31208.n142 a_34044_31208.t78 7.285
R134 a_34044_31208.n142 a_34044_31208.n141 14.37
R135 a_34044_31208.n141 a_34044_31208.t121 7.285
R136 a_34044_31208.n141 a_34044_31208.n140 14.37
R137 a_34044_31208.n140 a_34044_31208.t189 7.285
R138 a_34044_31208.n140 a_34044_31208.n139 14.395
R139 a_34044_31208.n139 a_34044_31208.t43 7.285
R140 a_34044_31208.n139 a_34044_31208.n138 14.37
R141 a_34044_31208.n138 a_34044_31208.t197 7.285
R142 a_34044_31208.n138 a_34044_31208.n137 14.37
R143 a_34044_31208.n137 a_34044_31208.t64 7.285
R144 a_34044_31208.n137 a_34044_31208.n136 14.37
R145 a_34044_31208.n136 a_34044_31208.t108 7.285
R146 a_34044_31208.n136 a_34044_31208.n135 15.728
R147 a_34044_31208.n135 a_34044_31208.t23 7.285
R148 a_34044_31208.n135 a_34044_31208.t90 21.655
R149 a_34044_31208.n134 a_34044_31208.n124 60.271
R150 a_34044_31208.n124 a_34044_31208.n133 7.74
R151 a_34044_31208.n133 a_34044_31208.t167 7.285
R152 a_34044_31208.n133 a_34044_31208.n132 14.37
R153 a_34044_31208.n132 a_34044_31208.t38 7.285
R154 a_34044_31208.n132 a_34044_31208.n131 14.37
R155 a_34044_31208.n131 a_34044_31208.t83 7.285
R156 a_34044_31208.n131 a_34044_31208.n130 14.37
R157 a_34044_31208.n130 a_34044_31208.t150 7.285
R158 a_34044_31208.n130 a_34044_31208.n129 14.395
R159 a_34044_31208.n129 a_34044_31208.t201 7.285
R160 a_34044_31208.n129 a_34044_31208.n128 14.37
R161 a_34044_31208.n128 a_34044_31208.t154 7.285
R162 a_34044_31208.n128 a_34044_31208.n127 14.37
R163 a_34044_31208.n127 a_34044_31208.t24 7.285
R164 a_34044_31208.n127 a_34044_31208.n126 14.37
R165 a_34044_31208.n126 a_34044_31208.t70 7.285
R166 a_34044_31208.n126 a_34044_31208.n125 15.728
R167 a_34044_31208.n125 a_34044_31208.t178 7.285
R168 a_34044_31208.n125 a_34044_31208.t50 21.655
R169 a_34044_31208.n124 a_34044_31208.n114 56.265
R170 a_34044_31208.n114 a_34044_31208.n123 7.74
R171 a_34044_31208.n123 a_34044_31208.t130 7.285
R172 a_34044_31208.n123 a_34044_31208.n122 14.37
R173 a_34044_31208.n122 a_34044_31208.t198 7.285
R174 a_34044_31208.n122 a_34044_31208.n121 14.37
R175 a_34044_31208.n121 a_34044_31208.t44 7.285
R176 a_34044_31208.n121 a_34044_31208.n120 14.37
R177 a_34044_31208.n120 a_34044_31208.t110 7.285
R178 a_34044_31208.n120 a_34044_31208.n119 14.395
R179 a_34044_31208.n119 a_34044_31208.t159 7.285
R180 a_34044_31208.n119 a_34044_31208.n118 14.37
R181 a_34044_31208.n118 a_34044_31208.t115 7.285
R182 a_34044_31208.n118 a_34044_31208.n117 14.37
R183 a_34044_31208.n117 a_34044_31208.t180 7.285
R184 a_34044_31208.n117 a_34044_31208.n116 14.37
R185 a_34044_31208.n116 a_34044_31208.t29 7.285
R186 a_34044_31208.n116 a_34044_31208.n115 15.728
R187 a_34044_31208.n115 a_34044_31208.t186 7.285
R188 a_34044_31208.n115 a_34044_31208.t58 21.655
R189 a_34044_31208.n114 a_34044_31208.n104 64.641
R190 a_34044_31208.n104 a_34044_31208.n113 7.74
R191 a_34044_31208.n113 a_34044_31208.t177 7.285
R192 a_34044_31208.n113 a_34044_31208.n112 14.37
R193 a_34044_31208.n112 a_34044_31208.t49 7.285
R194 a_34044_31208.n112 a_34044_31208.n111 14.37
R195 a_34044_31208.n111 a_34044_31208.t94 7.285
R196 a_34044_31208.n111 a_34044_31208.n110 14.37
R197 a_34044_31208.n110 a_34044_31208.t158 7.285
R198 a_34044_31208.n110 a_34044_31208.n109 14.395
R199 a_34044_31208.n109 a_34044_31208.t10 7.285
R200 a_34044_31208.n109 a_34044_31208.n108 14.37
R201 a_34044_31208.n108 a_34044_31208.t162 7.285
R202 a_34044_31208.n108 a_34044_31208.n107 14.37
R203 a_34044_31208.n107 a_34044_31208.t32 7.285
R204 a_34044_31208.n107 a_34044_31208.n106 14.37
R205 a_34044_31208.n106 a_34044_31208.t79 7.285
R206 a_34044_31208.n106 a_34044_31208.n105 15.728
R207 a_34044_31208.n105 a_34044_31208.t187 7.285
R208 a_34044_31208.n105 a_34044_31208.t59 21.655
R209 a_34044_31208.n104 a_34044_31208.n94 60.453
R210 a_34044_31208.n94 a_34044_31208.n103 7.74
R211 a_34044_31208.n103 a_34044_31208.t138 7.285
R212 a_34044_31208.n103 a_34044_31208.n102 14.37
R213 a_34044_31208.n102 a_34044_31208.t6 7.285
R214 a_34044_31208.n102 a_34044_31208.n101 14.37
R215 a_34044_31208.n101 a_34044_31208.t54 7.285
R216 a_34044_31208.n101 a_34044_31208.n100 14.37
R217 a_34044_31208.n100 a_34044_31208.t118 7.285
R218 a_34044_31208.n100 a_34044_31208.n99 14.395
R219 a_34044_31208.n99 a_34044_31208.t169 7.285
R220 a_34044_31208.n99 a_34044_31208.n98 14.37
R221 a_34044_31208.n98 a_34044_31208.t122 7.285
R222 a_34044_31208.n98 a_34044_31208.n97 14.37
R223 a_34044_31208.n97 a_34044_31208.t190 7.285
R224 a_34044_31208.n97 a_34044_31208.n96 14.37
R225 a_34044_31208.n96 a_34044_31208.t39 7.285
R226 a_34044_31208.n96 a_34044_31208.n95 15.728
R227 a_34044_31208.n95 a_34044_31208.t149 7.285
R228 a_34044_31208.n95 a_34044_31208.t20 21.655
R229 a_34044_31208.n94 a_34044_31208.n84 60.271
R230 a_34044_31208.n84 a_34044_31208.n93 7.74
R231 a_34044_31208.n93 a_34044_31208.t31 7.285
R232 a_34044_31208.n93 a_34044_31208.n92 14.37
R233 a_34044_31208.n92 a_34044_31208.t98 7.285
R234 a_34044_31208.n92 a_34044_31208.n91 14.37
R235 a_34044_31208.n91 a_34044_31208.t141 7.285
R236 a_34044_31208.n91 a_34044_31208.n90 14.37
R237 a_34044_31208.n90 a_34044_31208.t11 7.285
R238 a_34044_31208.n90 a_34044_31208.n89 14.395
R239 a_34044_31208.n89 a_34044_31208.t66 7.285
R240 a_34044_31208.n89 a_34044_31208.n88 14.37
R241 a_34044_31208.n88 a_34044_31208.t18 7.285
R242 a_34044_31208.n88 a_34044_31208.n87 14.37
R243 a_34044_31208.n87 a_34044_31208.t84 7.285
R244 a_34044_31208.n87 a_34044_31208.n86 14.37
R245 a_34044_31208.n86 a_34044_31208.t131 7.285
R246 a_34044_31208.n86 a_34044_31208.n85 15.728
R247 a_34044_31208.n85 a_34044_31208.t42 7.285
R248 a_34044_31208.n85 a_34044_31208.t109 21.655
R249 a_34044_31208.n84 a_34044_31208.n74 60.453
R250 a_34044_31208.n74 a_34044_31208.n83 7.74
R251 a_34044_31208.n83 a_34044_31208.t12 7.285
R252 a_34044_31208.n83 a_34044_31208.n82 14.37
R253 a_34044_31208.n82 a_34044_31208.t81 7.285
R254 a_34044_31208.n82 a_34044_31208.n81 14.37
R255 a_34044_31208.n81 a_34044_31208.t127 7.285
R256 a_34044_31208.n81 a_34044_31208.n80 14.37
R257 a_34044_31208.n80 a_34044_31208.t196 7.285
R258 a_34044_31208.n80 a_34044_31208.n79 14.395
R259 a_34044_31208.n79 a_34044_31208.t47 7.285
R260 a_34044_31208.n79 a_34044_31208.n78 14.37
R261 a_34044_31208.n78 a_34044_31208.t199 7.285
R262 a_34044_31208.n78 a_34044_31208.n77 14.37
R263 a_34044_31208.n77 a_34044_31208.t67 7.285
R264 a_34044_31208.n77 a_34044_31208.n76 14.37
R265 a_34044_31208.n76 a_34044_31208.t112 7.285
R266 a_34044_31208.n76 a_34044_31208.n75 15.728
R267 a_34044_31208.n75 a_34044_31208.t25 7.285
R268 a_34044_31208.n75 a_34044_31208.t91 21.655
R269 a_34044_31208.n74 a_34044_31208.n64 61
R270 a_34044_31208.n64 a_34044_31208.n73 7.74
R271 a_34044_31208.n73 a_34044_31208.t171 7.285
R272 a_34044_31208.n73 a_34044_31208.n72 14.37
R273 a_34044_31208.n72 a_34044_31208.t41 7.285
R274 a_34044_31208.n72 a_34044_31208.n71 14.37
R275 a_34044_31208.n71 a_34044_31208.t88 7.285
R276 a_34044_31208.n71 a_34044_31208.n70 14.37
R277 a_34044_31208.n70 a_34044_31208.t153 7.285
R278 a_34044_31208.n70 a_34044_31208.n69 14.395
R279 a_34044_31208.n69 a_34044_31208.t4 7.285
R280 a_34044_31208.n69 a_34044_31208.n68 14.37
R281 a_34044_31208.n68 a_34044_31208.t155 7.285
R282 a_34044_31208.n68 a_34044_31208.n67 14.37
R283 a_34044_31208.n67 a_34044_31208.t27 7.285
R284 a_34044_31208.n67 a_34044_31208.n66 14.37
R285 a_34044_31208.n66 a_34044_31208.t71 7.285
R286 a_34044_31208.n66 a_34044_31208.n65 15.728
R287 a_34044_31208.n65 a_34044_31208.t163 7.285
R288 a_34044_31208.n65 a_34044_31208.t33 21.655
R289 a_34044_31208.n64 a_34044_31208.n54 60.089
R290 a_34044_31208.n54 a_34044_31208.n63 7.74
R291 a_34044_31208.n63 a_34044_31208.t116 7.285
R292 a_34044_31208.n63 a_34044_31208.n62 14.37
R293 a_34044_31208.n62 a_34044_31208.t181 7.285
R294 a_34044_31208.n62 a_34044_31208.n61 14.37
R295 a_34044_31208.n61 a_34044_31208.t30 7.285
R296 a_34044_31208.n61 a_34044_31208.n60 14.37
R297 a_34044_31208.n60 a_34044_31208.t96 7.285
R298 a_34044_31208.n60 a_34044_31208.n59 14.395
R299 a_34044_31208.n59 a_34044_31208.t144 7.285
R300 a_34044_31208.n59 a_34044_31208.n58 14.37
R301 a_34044_31208.n58 a_34044_31208.t99 7.285
R302 a_34044_31208.n58 a_34044_31208.n57 14.37
R303 a_34044_31208.n57 a_34044_31208.t164 7.285
R304 a_34044_31208.n57 a_34044_31208.n56 14.37
R305 a_34044_31208.n56 a_34044_31208.t13 7.285
R306 a_34044_31208.n56 a_34044_31208.n55 15.728
R307 a_34044_31208.n55 a_34044_31208.t124 7.285
R308 a_34044_31208.n55 a_34044_31208.t191 21.655
R309 a_34044_31208.n54 a_34044_31208.n44 64.277
R310 a_34044_31208.n44 a_34044_31208.n53 7.74
R311 a_34044_31208.n53 a_34044_31208.t182 7.285
R312 a_34044_31208.n53 a_34044_31208.n52 14.37
R313 a_34044_31208.n52 a_34044_31208.t53 7.285
R314 a_34044_31208.n52 a_34044_31208.n51 14.37
R315 a_34044_31208.n51 a_34044_31208.t97 7.285
R316 a_34044_31208.n51 a_34044_31208.n50 14.37
R317 a_34044_31208.n50 a_34044_31208.t161 7.285
R318 a_34044_31208.n50 a_34044_31208.n49 14.395
R319 a_34044_31208.n49 a_34044_31208.t15 7.285
R320 a_34044_31208.n49 a_34044_31208.n48 14.37
R321 a_34044_31208.n48 a_34044_31208.t165 7.285
R322 a_34044_31208.n48 a_34044_31208.n47 14.37
R323 a_34044_31208.n47 a_34044_31208.t37 7.285
R324 a_34044_31208.n47 a_34044_31208.n46 14.37
R325 a_34044_31208.n46 a_34044_31208.t82 7.285
R326 a_34044_31208.n46 a_34044_31208.n45 15.728
R327 a_34044_31208.n45 a_34044_31208.t192 7.285
R328 a_34044_31208.n45 a_34044_31208.t62 21.655
R329 a_34044_31208.n44 a_34044_31208.n34 60.089
R330 a_34044_31208.n34 a_34044_31208.n43 7.74
R331 a_34044_31208.n43 a_34044_31208.t74 7.285
R332 a_34044_31208.n43 a_34044_31208.n42 14.37
R333 a_34044_31208.n42 a_34044_31208.t140 7.285
R334 a_34044_31208.n42 a_34044_31208.n41 14.37
R335 a_34044_31208.n41 a_34044_31208.t185 7.285
R336 a_34044_31208.n41 a_34044_31208.n40 14.37
R337 a_34044_31208.n40 a_34044_31208.t57 7.285
R338 a_34044_31208.n40 a_34044_31208.n39 14.395
R339 a_34044_31208.n39 a_34044_31208.t105 7.285
R340 a_34044_31208.n39 a_34044_31208.n38 14.37
R341 a_34044_31208.n38 a_34044_31208.t61 7.285
R342 a_34044_31208.n38 a_34044_31208.n37 14.37
R343 a_34044_31208.n37 a_34044_31208.t128 7.285
R344 a_34044_31208.n37 a_34044_31208.n36 14.37
R345 a_34044_31208.n36 a_34044_31208.t172 7.285
R346 a_34044_31208.n36 a_34044_31208.n35 15.728
R347 a_34044_31208.n35 a_34044_31208.t86 7.285
R348 a_34044_31208.n35 a_34044_31208.t152 21.655
R349 a_34044_31208.n34 a_34044_31208.n24 60.089
R350 a_34044_31208.n24 a_34044_31208.n33 7.74
R351 a_34044_31208.n33 a_34044_31208.t36 7.285
R352 a_34044_31208.n33 a_34044_31208.n32 14.37
R353 a_34044_31208.n32 a_34044_31208.t101 7.285
R354 a_34044_31208.n32 a_34044_31208.n31 14.37
R355 a_34044_31208.n31 a_34044_31208.t147 7.285
R356 a_34044_31208.n31 a_34044_31208.n30 14.37
R357 a_34044_31208.n30 a_34044_31208.t17 7.285
R358 a_34044_31208.n30 a_34044_31208.n29 14.395
R359 a_34044_31208.n29 a_34044_31208.t69 7.285
R360 a_34044_31208.n29 a_34044_31208.n28 14.37
R361 a_34044_31208.n28 a_34044_31208.t22 7.285
R362 a_34044_31208.n28 a_34044_31208.n27 14.37
R363 a_34044_31208.n27 a_34044_31208.t89 7.285
R364 a_34044_31208.n27 a_34044_31208.n26 14.37
R365 a_34044_31208.n26 a_34044_31208.t134 7.285
R366 a_34044_31208.n26 a_34044_31208.n25 15.728
R367 a_34044_31208.n25 a_34044_31208.t46 7.285
R368 a_34044_31208.n25 a_34044_31208.t114 21.655
R369 a_34044_31208.n24 a_34044_31208.n23 67.83
R370 a_34044_31208.n23 a_34044_31208.t148 7.285
R371 a_34044_31208.n23 a_34044_31208.n22 14.37
R372 a_34044_31208.n22 a_34044_31208.t19 7.285
R373 a_34044_31208.n22 a_34044_31208.n21 14.37
R374 a_34044_31208.n21 a_34044_31208.t65 7.285
R375 a_34044_31208.n21 a_34044_31208.n20 14.37
R376 a_34044_31208.n20 a_34044_31208.t132 7.285
R377 a_34044_31208.n20 a_34044_31208.n19 14.395
R378 a_34044_31208.n19 a_34044_31208.t179 7.285
R379 a_34044_31208.n19 a_34044_31208.n18 14.37
R380 a_34044_31208.n18 a_34044_31208.t135 7.285
R381 a_34044_31208.n18 a_34044_31208.n17 14.37
R382 a_34044_31208.n17 a_34044_31208.t200 7.285
R383 a_34044_31208.n17 a_34044_31208.n16 14.37
R384 a_34044_31208.n16 a_34044_31208.t51 7.285
R385 a_34044_31208.n16 a_34044_31208.n15 15.728
R386 a_34044_31208.n15 a_34044_31208.t8 7.285
R387 a_34044_31208.n15 a_34044_31208.t76 21.655
R388 a_34044_31208.n12 a_34044_31208.t168 21.738
R389 a_34044_31208.n12 a_34044_31208.t102 7.262
R390 a_34044_31208.n11 a_34044_31208.t188 7.262
R391 a_34044_31208.n11 a_34044_31208.n12 15.847
R392 a_34044_31208.n10 a_34044_31208.t142 7.262
R393 a_34044_31208.n10 a_34044_31208.n11 14.475
R394 a_34044_31208.n8 a_34044_31208.t77 21.087
R395 a_34044_31208.n7 a_34044_31208.t123 7.262
R396 a_34044_31208.n7 a_34044_31208.n8 7.911
R397 a_34044_31208.n6 a_34044_31208.t72 7.262
R398 a_34044_31208.n6 a_34044_31208.n7 14.5
R399 a_34044_31208.n5 a_34044_31208.t5 7.262
R400 a_34044_31208.n5 a_34044_31208.n6 14.475
R401 a_34044_31208.n4 a_34044_31208.t157 7.262
R402 a_34044_31208.n4 a_34044_31208.n5 14.475
R403 a_34044_31208.n3 a_34044_31208.t93 7.262
R404 a_34044_31208.n3 a_34044_31208.n4 14.475
R405 a_34044_31208.n204 a_34044_31208.n1 3.542
R406 a_34044_31208.n1 a_34044_31208.t2 19.8
R407 a_34044_31208.n1 a_34044_31208.t0 19.8
R408 a_66167_26022.n3 a_66167_26022.t4 389.181
R409 a_66167_26022.n0 a_66167_26022.t5 256.987
R410 a_66167_26022.n2 a_66167_26022.t3 212.079
R411 a_66167_26022.n3 a_66167_26022.t7 174.888
R412 a_66167_26022.n0 a_66167_26022.t8 163.801
R413 a_66167_26022.n6 a_66167_26022.n5 161.578
R414 a_66167_26022.n1 a_66167_26022.t6 139.779
R415 a_66167_26022.n1 a_66167_26022.n0 129.263
R416 a_66167_26022.n4 a_66167_26022.n3 102.015
R417 a_66167_26022.n6 a_66167_26022.t2 63.321
R418 a_66167_26022.t0 a_66167_26022.n6 63.321
R419 a_66167_26022.n4 a_66167_26022.t1 46.071
R420 a_66167_26022.n5 a_66167_26022.n2 37.442
R421 a_66167_26022.n5 a_66167_26022.n4 23.54
R422 a_66167_26022.n2 a_66167_26022.n1 22.639
R423 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.n2 1158.04
R424 Fvco_By4_QPH_bar.t8 Fvco_By4_QPH_bar.t7 731.89
R425 Fvco_By4_QPH_bar.t3 Fvco_By4_QPH_bar.t12 719.978
R426 Fvco_By4_QPH_bar.t6 Fvco_By4_QPH_bar.t16 710.965
R427 Fvco_By4_QPH_bar.t5 Fvco_By4_QPH_bar.t17 710.965
R428 Fvco_By4_QPH_bar.t4 Fvco_By4_QPH_bar.t11 710.965
R429 Fvco_By4_QPH_bar.t16 Fvco_By4_QPH_bar.t15 579.889
R430 Fvco_By4_QPH_bar.t17 Fvco_By4_QPH_bar.t13 579.889
R431 Fvco_By4_QPH_bar.t11 Fvco_By4_QPH_bar.t10 579.889
R432 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.t5 570.03
R433 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.t4 563.963
R434 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t6 557.83
R435 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n0 458.189
R436 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.n5 435.858
R437 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t14 417.917
R438 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.t9 414.213
R439 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.t2 414.167
R440 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.t3 245.573
R441 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.t8 244.389
R442 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n7 188.615
R443 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n4 149.023
R444 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.n6 130.017
R445 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t0 69.215
R446 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n1 50.411
R447 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t1 39.949
R448 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.n3 1.452
R449 a_26368_16652.t24 a_26368_16652.t49 1273.78
R450 a_26368_16652.n0 a_26368_16652.t24 182.777
R451 a_26368_16652.n0 a_26368_16652.t0 127.728
R452 a_26368_16652.t24 a_26368_16652.t52 127.098
R453 a_26368_16652.t24 a_26368_16652.t21 113.753
R454 a_26368_16652.t24 a_26368_16652.t27 113.753
R455 a_26368_16652.t24 a_26368_16652.t42 113.753
R456 a_26368_16652.t24 a_26368_16652.t57 113.753
R457 a_26368_16652.t24 a_26368_16652.t51 113.753
R458 a_26368_16652.t24 a_26368_16652.t3 113.753
R459 a_26368_16652.t24 a_26368_16652.t16 113.753
R460 a_26368_16652.t24 a_26368_16652.t32 113.753
R461 a_26368_16652.t24 a_26368_16652.t28 113.753
R462 a_26368_16652.t24 a_26368_16652.t41 113.753
R463 a_26368_16652.t24 a_26368_16652.t56 113.753
R464 a_26368_16652.t24 a_26368_16652.t12 113.753
R465 a_26368_16652.t24 a_26368_16652.t35 113.753
R466 a_26368_16652.t24 a_26368_16652.t47 113.753
R467 a_26368_16652.t24 a_26368_16652.t6 113.753
R468 a_26368_16652.t24 a_26368_16652.t59 113.753
R469 a_26368_16652.t24 a_26368_16652.t13 113.753
R470 a_26368_16652.t24 a_26368_16652.t29 113.753
R471 a_26368_16652.t24 a_26368_16652.t43 113.753
R472 a_26368_16652.t24 a_26368_16652.t22 113.753
R473 a_26368_16652.t24 a_26368_16652.t8 113.753
R474 a_26368_16652.t24 a_26368_16652.t19 113.753
R475 a_26368_16652.t24 a_26368_16652.t37 113.753
R476 a_26368_16652.t24 a_26368_16652.t33 113.753
R477 a_26368_16652.t24 a_26368_16652.t45 113.753
R478 a_26368_16652.t24 a_26368_16652.t4 113.753
R479 a_26368_16652.t24 a_26368_16652.t17 113.753
R480 a_26368_16652.t24 a_26368_16652.t36 113.753
R481 a_26368_16652.t24 a_26368_16652.t48 113.753
R482 a_26368_16652.t24 a_26368_16652.t7 113.753
R483 a_26368_16652.t24 a_26368_16652.t2 113.753
R484 a_26368_16652.t24 a_26368_16652.t14 113.753
R485 a_26368_16652.t24 a_26368_16652.t30 113.753
R486 a_26368_16652.t24 a_26368_16652.t44 113.753
R487 a_26368_16652.t24 a_26368_16652.t23 113.753
R488 a_26368_16652.t24 a_26368_16652.t53 113.753
R489 a_26368_16652.t24 a_26368_16652.t9 113.753
R490 a_26368_16652.t24 a_26368_16652.t20 113.753
R491 a_26368_16652.t24 a_26368_16652.t38 113.753
R492 a_26368_16652.t24 a_26368_16652.t34 113.753
R493 a_26368_16652.t24 a_26368_16652.t46 113.753
R494 a_26368_16652.t24 a_26368_16652.t5 113.753
R495 a_26368_16652.t24 a_26368_16652.t18 113.753
R496 a_26368_16652.t24 a_26368_16652.t50 113.753
R497 a_26368_16652.t24 a_26368_16652.t58 113.753
R498 a_26368_16652.t24 a_26368_16652.t15 113.753
R499 a_26368_16652.t24 a_26368_16652.t31 113.753
R500 a_26368_16652.t24 a_26368_16652.t26 113.753
R501 a_26368_16652.t24 a_26368_16652.t40 113.753
R502 a_26368_16652.t24 a_26368_16652.t55 113.753
R503 a_26368_16652.t24 a_26368_16652.t11 113.753
R504 a_26368_16652.t24 a_26368_16652.t54 113.753
R505 a_26368_16652.t24 a_26368_16652.t10 113.753
R506 a_26368_16652.t24 a_26368_16652.t25 113.753
R507 a_26368_16652.t24 a_26368_16652.t39 113.753
R508 a_26368_16652.t1 a_26368_16652.n0 57.482
R509 a_28736_17218.n0 a_28736_17218.n3 75.71
R510 a_28736_17218.n4 a_28736_17218.n5 75.708
R511 a_28736_17218.n2 a_28736_17218.n1 75.707
R512 a_28736_17218.n3 a_28736_17218.n2 75.707
R513 a_28736_17218.n1 a_28736_17218.n6 75.707
R514 a_28736_17218.n0 a_28736_17218.n4 75.706
R515 a_28736_17218.n0 a_28736_17218.t11 17.401
R516 a_28736_17218.n4 a_28736_17218.t7 17.401
R517 a_28736_17218.n3 a_28736_17218.t3 17.401
R518 a_28736_17218.n2 a_28736_17218.t8 17.401
R519 a_28736_17218.n1 a_28736_17218.t9 17.401
R520 a_28736_17218.n5 a_28736_17218.t10 17.4
R521 a_28736_17218.n5 a_28736_17218.t6 17.4
R522 a_28736_17218.n4 a_28736_17218.t13 17.4
R523 a_28736_17218.n3 a_28736_17218.t2 17.4
R524 a_28736_17218.n2 a_28736_17218.t1 17.4
R525 a_28736_17218.n1 a_28736_17218.t12 17.4
R526 a_28736_17218.n6 a_28736_17218.t4 17.4
R527 a_28736_17218.n6 a_28736_17218.t5 17.4
R528 a_28736_17218.t0 a_28736_17218.n0 17.4
R529 a_28994_17218.n0 a_28994_17218.n4 75.71
R530 a_28994_17218.n2 a_28994_17218.n1 75.707
R531 a_28994_17218.n3 a_28994_17218.n2 75.707
R532 a_28994_17218.n4 a_28994_17218.n3 75.707
R533 a_28994_17218.n1 a_28994_17218.n6 75.707
R534 a_28994_17218.n0 a_28994_17218.n5 75.707
R535 a_28994_17218.n0 a_28994_17218.t11 17.401
R536 a_28994_17218.n4 a_28994_17218.t10 17.401
R537 a_28994_17218.n3 a_28994_17218.t12 17.401
R538 a_28994_17218.n2 a_28994_17218.t7 17.401
R539 a_28994_17218.n1 a_28994_17218.t8 17.401
R540 a_28994_17218.n5 a_28994_17218.t9 17.4
R541 a_28994_17218.n5 a_28994_17218.t2 17.4
R542 a_28994_17218.n4 a_28994_17218.t3 17.4
R543 a_28994_17218.n3 a_28994_17218.t0 17.4
R544 a_28994_17218.n2 a_28994_17218.t4 17.4
R545 a_28994_17218.n1 a_28994_17218.t5 17.4
R546 a_28994_17218.n6 a_28994_17218.t13 17.4
R547 a_28994_17218.n6 a_28994_17218.t1 17.4
R548 a_28994_17218.t6 a_28994_17218.n0 17.4
R549 a_23414_5032.t2 a_23414_5032.t41 1273.78
R550 a_23414_5032.t2 a_23414_5032.t14 345.988
R551 a_23414_5032.t14 a_23414_5032.t49 126.864
R552 a_23414_5032.t14 a_23414_5032.t5 113.753
R553 a_23414_5032.t14 a_23414_5032.t3 113.753
R554 a_23414_5032.t14 a_23414_5032.t15 113.753
R555 a_23414_5032.t14 a_23414_5032.t37 113.753
R556 a_23414_5032.t14 a_23414_5032.t33 113.753
R557 a_23414_5032.t14 a_23414_5032.t31 113.753
R558 a_23414_5032.t14 a_23414_5032.t30 113.753
R559 a_23414_5032.t14 a_23414_5032.t7 113.753
R560 a_23414_5032.t14 a_23414_5032.t39 113.753
R561 a_23414_5032.t14 a_23414_5032.t36 113.753
R562 a_23414_5032.t14 a_23414_5032.t34 113.753
R563 a_23414_5032.t14 a_23414_5032.t45 113.753
R564 a_23414_5032.t14 a_23414_5032.t11 113.753
R565 a_23414_5032.t14 a_23414_5032.t8 113.753
R566 a_23414_5032.t14 a_23414_5032.t6 113.753
R567 a_23414_5032.t14 a_23414_5032.t4 113.753
R568 a_23414_5032.t14 a_23414_5032.t21 113.753
R569 a_23414_5032.t14 a_23414_5032.t17 113.753
R570 a_23414_5032.t14 a_23414_5032.t35 113.753
R571 a_23414_5032.t14 a_23414_5032.t56 113.753
R572 a_23414_5032.t14 a_23414_5032.t51 113.753
R573 a_23414_5032.t14 a_23414_5032.t47 113.753
R574 a_23414_5032.t14 a_23414_5032.t24 113.753
R575 a_23414_5032.t14 a_23414_5032.t58 113.753
R576 a_23414_5032.t14 a_23414_5032.t55 113.753
R577 a_23414_5032.t14 a_23414_5032.t52 113.753
R578 a_23414_5032.t14 a_23414_5032.t9 113.753
R579 a_23414_5032.t14 a_23414_5032.t28 113.753
R580 a_23414_5032.t14 a_23414_5032.t25 113.753
R581 a_23414_5032.t14 a_23414_5032.t23 113.753
R582 a_23414_5032.t14 a_23414_5032.t20 113.753
R583 a_23414_5032.t14 a_23414_5032.t27 113.753
R584 a_23414_5032.t14 a_23414_5032.t26 113.753
R585 a_23414_5032.t14 a_23414_5032.t42 113.753
R586 a_23414_5032.t14 a_23414_5032.t60 113.753
R587 a_23414_5032.t14 a_23414_5032.t59 113.753
R588 a_23414_5032.t14 a_23414_5032.t57 113.753
R589 a_23414_5032.t14 a_23414_5032.t54 113.753
R590 a_23414_5032.t14 a_23414_5032.t29 113.753
R591 a_23414_5032.t14 a_23414_5032.t13 113.753
R592 a_23414_5032.t14 a_23414_5032.t12 113.753
R593 a_23414_5032.t14 a_23414_5032.t10 113.753
R594 a_23414_5032.t14 a_23414_5032.t18 113.753
R595 a_23414_5032.t14 a_23414_5032.t44 113.753
R596 a_23414_5032.t14 a_23414_5032.t43 113.753
R597 a_23414_5032.t14 a_23414_5032.t40 113.753
R598 a_23414_5032.t14 a_23414_5032.t38 113.753
R599 a_23414_5032.t14 a_23414_5032.t22 113.753
R600 a_23414_5032.t14 a_23414_5032.t19 113.753
R601 a_23414_5032.t14 a_23414_5032.t16 113.753
R602 a_23414_5032.t14 a_23414_5032.t32 113.753
R603 a_23414_5032.t14 a_23414_5032.t53 113.753
R604 a_23414_5032.t14 a_23414_5032.t50 113.753
R605 a_23414_5032.t14 a_23414_5032.t48 113.753
R606 a_23414_5032.t14 a_23414_5032.t46 113.753
R607 a_23414_5032.t0 a_23414_5032.t2 82.513
R608 a_23414_5032.t2 a_23414_5032.t1 34.838
R609 a_26690_784.n1 a_26690_784.t2 434.481
R610 a_26690_784.n0 a_26690_784.t3 217.163
R611 a_26690_784.t1 a_26690_784.n1 52.152
R612 a_26690_784.n0 a_26690_784.t0 3.106
R613 a_26690_784.n1 a_26690_784.n0 0.879
R614 a_1026_45630.n0 a_1026_45630.t2 16.252
R615 a_1026_45630.t0 a_1026_45630.n0 16.252
R616 a_1026_45630.n0 a_1026_45630.n1 1.568
R617 a_1026_45630.n1 a_1026_45630.n201 2.477
R618 a_1026_45630.n201 a_1026_45630.t3 19.8
R619 a_1026_45630.n201 a_1026_45630.t1 19.8
R620 a_1026_45630.n1 a_1026_45630.n200 133.854
R621 a_1026_45630.n200 a_1026_45630.n190 206.115
R622 a_1026_45630.n190 a_1026_45630.n199 7.345
R623 a_1026_45630.n199 a_1026_45630.t187 7.285
R624 a_1026_45630.n199 a_1026_45630.n198 14.37
R625 a_1026_45630.n198 a_1026_45630.t54 7.285
R626 a_1026_45630.n198 a_1026_45630.n197 14.37
R627 a_1026_45630.n197 a_1026_45630.t104 7.285
R628 a_1026_45630.n197 a_1026_45630.n196 14.37
R629 a_1026_45630.n196 a_1026_45630.t169 7.285
R630 a_1026_45630.n196 a_1026_45630.n195 14.395
R631 a_1026_45630.n195 a_1026_45630.t23 7.285
R632 a_1026_45630.n195 a_1026_45630.n194 14.37
R633 a_1026_45630.n194 a_1026_45630.t176 7.285
R634 a_1026_45630.n194 a_1026_45630.n193 14.37
R635 a_1026_45630.n193 a_1026_45630.t40 7.285
R636 a_1026_45630.n193 a_1026_45630.n192 14.37
R637 a_1026_45630.n192 a_1026_45630.t93 7.285
R638 a_1026_45630.n192 a_1026_45630.n191 15.728
R639 a_1026_45630.n191 a_1026_45630.t199 7.285
R640 a_1026_45630.n191 a_1026_45630.t66 21.655
R641 a_1026_45630.n190 a_1026_45630.n180 213.178
R642 a_1026_45630.n180 a_1026_45630.n189 7.345
R643 a_1026_45630.n189 a_1026_45630.t186 7.285
R644 a_1026_45630.n189 a_1026_45630.n188 14.37
R645 a_1026_45630.n188 a_1026_45630.t53 7.285
R646 a_1026_45630.n188 a_1026_45630.n187 14.37
R647 a_1026_45630.n187 a_1026_45630.t103 7.285
R648 a_1026_45630.n187 a_1026_45630.n186 14.37
R649 a_1026_45630.n186 a_1026_45630.t168 7.285
R650 a_1026_45630.n186 a_1026_45630.n185 14.395
R651 a_1026_45630.n185 a_1026_45630.t22 7.285
R652 a_1026_45630.n185 a_1026_45630.n184 14.37
R653 a_1026_45630.n184 a_1026_45630.t175 7.285
R654 a_1026_45630.n184 a_1026_45630.n183 14.37
R655 a_1026_45630.n183 a_1026_45630.t39 7.285
R656 a_1026_45630.n183 a_1026_45630.n182 14.37
R657 a_1026_45630.n182 a_1026_45630.t92 7.285
R658 a_1026_45630.n182 a_1026_45630.n181 15.728
R659 a_1026_45630.n181 a_1026_45630.t198 7.285
R660 a_1026_45630.n181 a_1026_45630.t65 21.655
R661 a_1026_45630.n180 a_1026_45630.n170 220.884
R662 a_1026_45630.n170 a_1026_45630.n179 7.345
R663 a_1026_45630.n179 a_1026_45630.t27 7.285
R664 a_1026_45630.n179 a_1026_45630.n178 14.37
R665 a_1026_45630.n178 a_1026_45630.t97 7.285
R666 a_1026_45630.n178 a_1026_45630.n177 14.37
R667 a_1026_45630.n177 a_1026_45630.t140 7.285
R668 a_1026_45630.n177 a_1026_45630.n176 14.37
R669 a_1026_45630.n176 a_1026_45630.t10 7.285
R670 a_1026_45630.n176 a_1026_45630.n175 14.395
R671 a_1026_45630.n175 a_1026_45630.t57 7.285
R672 a_1026_45630.n175 a_1026_45630.n174 14.37
R673 a_1026_45630.n174 a_1026_45630.t14 7.285
R674 a_1026_45630.n174 a_1026_45630.n173 14.37
R675 a_1026_45630.n173 a_1026_45630.t80 7.285
R676 a_1026_45630.n173 a_1026_45630.n172 14.37
R677 a_1026_45630.n172 a_1026_45630.t126 7.285
R678 a_1026_45630.n172 a_1026_45630.n171 15.728
R679 a_1026_45630.n171 a_1026_45630.t38 7.285
R680 a_1026_45630.n171 a_1026_45630.t110 21.655
R681 a_1026_45630.n170 a_1026_45630.n160 206.115
R682 a_1026_45630.n160 a_1026_45630.n169 7.345
R683 a_1026_45630.n169 a_1026_45630.t69 7.285
R684 a_1026_45630.n169 a_1026_45630.n168 14.37
R685 a_1026_45630.n168 a_1026_45630.t137 7.285
R686 a_1026_45630.n168 a_1026_45630.n167 14.37
R687 a_1026_45630.n167 a_1026_45630.t183 7.285
R688 a_1026_45630.n167 a_1026_45630.n166 14.37
R689 a_1026_45630.n166 a_1026_45630.t47 7.285
R690 a_1026_45630.n166 a_1026_45630.n165 14.395
R691 a_1026_45630.n165 a_1026_45630.t100 7.285
R692 a_1026_45630.n165 a_1026_45630.n164 14.37
R693 a_1026_45630.n164 a_1026_45630.t52 7.285
R694 a_1026_45630.n164 a_1026_45630.n163 14.37
R695 a_1026_45630.n163 a_1026_45630.t120 7.285
R696 a_1026_45630.n163 a_1026_45630.n162 14.37
R697 a_1026_45630.n162 a_1026_45630.t166 7.285
R698 a_1026_45630.n162 a_1026_45630.n161 15.728
R699 a_1026_45630.n161 a_1026_45630.t78 7.285
R700 a_1026_45630.n161 a_1026_45630.t145 21.655
R701 a_1026_45630.n160 a_1026_45630.n150 227.947
R702 a_1026_45630.n150 a_1026_45630.n159 7.345
R703 a_1026_45630.n159 a_1026_45630.t106 7.285
R704 a_1026_45630.n159 a_1026_45630.n158 14.37
R705 a_1026_45630.n158 a_1026_45630.t174 7.285
R706 a_1026_45630.n158 a_1026_45630.n157 14.37
R707 a_1026_45630.n157 a_1026_45630.t20 7.285
R708 a_1026_45630.n157 a_1026_45630.n156 14.37
R709 a_1026_45630.n156 a_1026_45630.t88 7.285
R710 a_1026_45630.n156 a_1026_45630.n155 14.395
R711 a_1026_45630.n155 a_1026_45630.t136 7.285
R712 a_1026_45630.n155 a_1026_45630.n154 14.37
R713 a_1026_45630.n154 a_1026_45630.t94 7.285
R714 a_1026_45630.n154 a_1026_45630.n153 14.37
R715 a_1026_45630.n153 a_1026_45630.t158 7.285
R716 a_1026_45630.n153 a_1026_45630.n152 14.37
R717 a_1026_45630.n152 a_1026_45630.t203 7.285
R718 a_1026_45630.n152 a_1026_45630.n151 15.728
R719 a_1026_45630.n151 a_1026_45630.t162 7.285
R720 a_1026_45630.n151 a_1026_45630.t29 21.655
R721 a_1026_45630.n150 a_1026_45630.n140 221.526
R722 a_1026_45630.n140 a_1026_45630.n149 7.345
R723 a_1026_45630.n149 a_1026_45630.t142 7.285
R724 a_1026_45630.n149 a_1026_45630.n148 14.37
R725 a_1026_45630.n148 a_1026_45630.t13 7.285
R726 a_1026_45630.n148 a_1026_45630.n147 14.37
R727 a_1026_45630.n147 a_1026_45630.t55 7.285
R728 a_1026_45630.n147 a_1026_45630.n146 14.37
R729 a_1026_45630.n146 a_1026_45630.t125 7.285
R730 a_1026_45630.n146 a_1026_45630.n145 14.395
R731 a_1026_45630.n145 a_1026_45630.t178 7.285
R732 a_1026_45630.n145 a_1026_45630.n144 14.37
R733 a_1026_45630.n144 a_1026_45630.t130 7.285
R734 a_1026_45630.n144 a_1026_45630.n143 14.37
R735 a_1026_45630.n143 a_1026_45630.t197 7.285
R736 a_1026_45630.n143 a_1026_45630.n142 14.37
R737 a_1026_45630.n142 a_1026_45630.t42 7.285
R738 a_1026_45630.n142 a_1026_45630.n141 15.728
R739 a_1026_45630.n141 a_1026_45630.t156 7.285
R740 a_1026_45630.n141 a_1026_45630.t25 21.655
R741 a_1026_45630.n140 a_1026_45630.n130 206.115
R742 a_1026_45630.n130 a_1026_45630.n139 7.345
R743 a_1026_45630.n139 a_1026_45630.t51 7.285
R744 a_1026_45630.n139 a_1026_45630.n138 14.37
R745 a_1026_45630.n138 a_1026_45630.t119 7.285
R746 a_1026_45630.n138 a_1026_45630.n137 14.37
R747 a_1026_45630.n137 a_1026_45630.t165 7.285
R748 a_1026_45630.n137 a_1026_45630.n136 14.37
R749 a_1026_45630.n136 a_1026_45630.t31 7.285
R750 a_1026_45630.n136 a_1026_45630.n135 14.395
R751 a_1026_45630.n135 a_1026_45630.t86 7.285
R752 a_1026_45630.n135 a_1026_45630.n134 14.37
R753 a_1026_45630.n134 a_1026_45630.t36 7.285
R754 a_1026_45630.n134 a_1026_45630.n133 14.37
R755 a_1026_45630.n133 a_1026_45630.t108 7.285
R756 a_1026_45630.n133 a_1026_45630.n132 14.37
R757 a_1026_45630.n132 a_1026_45630.t152 7.285
R758 a_1026_45630.n132 a_1026_45630.n131 15.728
R759 a_1026_45630.n131 a_1026_45630.t62 7.285
R760 a_1026_45630.n131 a_1026_45630.t132 21.655
R761 a_1026_45630.n130 a_1026_45630.n120 213.178
R762 a_1026_45630.n120 a_1026_45630.n129 7.345
R763 a_1026_45630.n129 a_1026_45630.t185 7.285
R764 a_1026_45630.n129 a_1026_45630.n128 14.37
R765 a_1026_45630.n128 a_1026_45630.t50 7.285
R766 a_1026_45630.n128 a_1026_45630.n127 14.37
R767 a_1026_45630.n127 a_1026_45630.t99 7.285
R768 a_1026_45630.n127 a_1026_45630.n126 14.37
R769 a_1026_45630.n126 a_1026_45630.t164 7.285
R770 a_1026_45630.n126 a_1026_45630.n125 14.395
R771 a_1026_45630.n125 a_1026_45630.t19 7.285
R772 a_1026_45630.n125 a_1026_45630.n124 14.37
R773 a_1026_45630.n124 a_1026_45630.t171 7.285
R774 a_1026_45630.n124 a_1026_45630.n123 14.37
R775 a_1026_45630.n123 a_1026_45630.t35 7.285
R776 a_1026_45630.n123 a_1026_45630.n122 14.37
R777 a_1026_45630.n122 a_1026_45630.t84 7.285
R778 a_1026_45630.n122 a_1026_45630.n121 15.728
R779 a_1026_45630.n121 a_1026_45630.t194 7.285
R780 a_1026_45630.n121 a_1026_45630.t61 21.655
R781 a_1026_45630.n120 a_1026_45630.n119 279.829
R782 a_1026_45630.n119 a_1026_45630.n109 183.395
R783 a_1026_45630.n109 a_1026_45630.n118 7.345
R784 a_1026_45630.n118 a_1026_45630.t83 7.285
R785 a_1026_45630.n118 a_1026_45630.n117 14.37
R786 a_1026_45630.n117 a_1026_45630.t151 7.285
R787 a_1026_45630.n117 a_1026_45630.n116 14.37
R788 a_1026_45630.n116 a_1026_45630.t196 7.285
R789 a_1026_45630.n116 a_1026_45630.n115 14.37
R790 a_1026_45630.n115 a_1026_45630.t63 7.285
R791 a_1026_45630.n115 a_1026_45630.n114 14.395
R792 a_1026_45630.n114 a_1026_45630.t114 7.285
R793 a_1026_45630.n114 a_1026_45630.n113 14.37
R794 a_1026_45630.n113 a_1026_45630.t68 7.285
R795 a_1026_45630.n113 a_1026_45630.n112 14.37
R796 a_1026_45630.n112 a_1026_45630.t135 7.285
R797 a_1026_45630.n112 a_1026_45630.n111 14.37
R798 a_1026_45630.n111 a_1026_45630.t181 7.285
R799 a_1026_45630.n111 a_1026_45630.n110 15.728
R800 a_1026_45630.n110 a_1026_45630.t141 7.285
R801 a_1026_45630.n110 a_1026_45630.t11 21.655
R802 a_1026_45630.n109 a_1026_45630.n99 228.589
R803 a_1026_45630.n99 a_1026_45630.n108 7.345
R804 a_1026_45630.n108 a_1026_45630.t101 7.285
R805 a_1026_45630.n108 a_1026_45630.n107 14.37
R806 a_1026_45630.n107 a_1026_45630.t167 7.285
R807 a_1026_45630.n107 a_1026_45630.n106 14.37
R808 a_1026_45630.n106 a_1026_45630.t16 7.285
R809 a_1026_45630.n106 a_1026_45630.n105 14.37
R810 a_1026_45630.n105 a_1026_45630.t82 7.285
R811 a_1026_45630.n105 a_1026_45630.n104 14.395
R812 a_1026_45630.n104 a_1026_45630.t134 7.285
R813 a_1026_45630.n104 a_1026_45630.n103 14.37
R814 a_1026_45630.n103 a_1026_45630.t90 7.285
R815 a_1026_45630.n103 a_1026_45630.n102 14.37
R816 a_1026_45630.n102 a_1026_45630.t154 7.285
R817 a_1026_45630.n102 a_1026_45630.n101 14.37
R818 a_1026_45630.n101 a_1026_45630.t200 7.285
R819 a_1026_45630.n101 a_1026_45630.n100 15.728
R820 a_1026_45630.n100 a_1026_45630.t113 7.285
R821 a_1026_45630.n100 a_1026_45630.t179 21.655
R822 a_1026_45630.n99 a_1026_45630.n89 213.178
R823 a_1026_45630.n89 a_1026_45630.n98 7.345
R824 a_1026_45630.n98 a_1026_45630.t9 7.285
R825 a_1026_45630.n98 a_1026_45630.n97 14.37
R826 a_1026_45630.n97 a_1026_45630.t74 7.285
R827 a_1026_45630.n97 a_1026_45630.n96 14.37
R828 a_1026_45630.n96 a_1026_45630.t122 7.285
R829 a_1026_45630.n96 a_1026_45630.n95 14.37
R830 a_1026_45630.n95 a_1026_45630.t189 7.285
R831 a_1026_45630.n95 a_1026_45630.n94 14.395
R832 a_1026_45630.n94 a_1026_45630.t41 7.285
R833 a_1026_45630.n94 a_1026_45630.n93 14.37
R834 a_1026_45630.n93 a_1026_45630.t192 7.285
R835 a_1026_45630.n93 a_1026_45630.n92 14.37
R836 a_1026_45630.n92 a_1026_45630.t58 7.285
R837 a_1026_45630.n92 a_1026_45630.n91 14.37
R838 a_1026_45630.n91 a_1026_45630.t111 7.285
R839 a_1026_45630.n91 a_1026_45630.n90 15.728
R840 a_1026_45630.n90 a_1026_45630.t21 7.285
R841 a_1026_45630.n90 a_1026_45630.t91 21.655
R842 a_1026_45630.n89 a_1026_45630.n79 206.115
R843 a_1026_45630.n79 a_1026_45630.n88 7.345
R844 a_1026_45630.n88 a_1026_45630.t46 7.285
R845 a_1026_45630.n88 a_1026_45630.n87 14.37
R846 a_1026_45630.n87 a_1026_45630.t115 7.285
R847 a_1026_45630.n87 a_1026_45630.n86 14.37
R848 a_1026_45630.n86 a_1026_45630.t160 7.285
R849 a_1026_45630.n86 a_1026_45630.n85 14.37
R850 a_1026_45630.n85 a_1026_45630.t28 7.285
R851 a_1026_45630.n85 a_1026_45630.n84 14.395
R852 a_1026_45630.n84 a_1026_45630.t81 7.285
R853 a_1026_45630.n84 a_1026_45630.n83 14.37
R854 a_1026_45630.n83 a_1026_45630.t32 7.285
R855 a_1026_45630.n83 a_1026_45630.n82 14.37
R856 a_1026_45630.n82 a_1026_45630.t102 7.285
R857 a_1026_45630.n82 a_1026_45630.n81 14.37
R858 a_1026_45630.n81 a_1026_45630.t146 7.285
R859 a_1026_45630.n81 a_1026_45630.n80 15.728
R860 a_1026_45630.n80 a_1026_45630.t56 7.285
R861 a_1026_45630.n80 a_1026_45630.t127 21.655
R862 a_1026_45630.n79 a_1026_45630.n69 213.178
R863 a_1026_45630.n69 a_1026_45630.n78 7.345
R864 a_1026_45630.n78 a_1026_45630.t98 7.285
R865 a_1026_45630.n78 a_1026_45630.n77 14.37
R866 a_1026_45630.n77 a_1026_45630.t161 7.285
R867 a_1026_45630.n77 a_1026_45630.n76 14.37
R868 a_1026_45630.n76 a_1026_45630.t8 7.285
R869 a_1026_45630.n76 a_1026_45630.n75 14.37
R870 a_1026_45630.n75 a_1026_45630.t75 7.285
R871 a_1026_45630.n75 a_1026_45630.n74 14.395
R872 a_1026_45630.n74 a_1026_45630.t128 7.285
R873 a_1026_45630.n74 a_1026_45630.n73 14.37
R874 a_1026_45630.n73 a_1026_45630.t79 7.285
R875 a_1026_45630.n73 a_1026_45630.n72 14.37
R876 a_1026_45630.n72 a_1026_45630.t149 7.285
R877 a_1026_45630.n72 a_1026_45630.n71 14.37
R878 a_1026_45630.n71 a_1026_45630.t193 7.285
R879 a_1026_45630.n71 a_1026_45630.n70 15.728
R880 a_1026_45630.n70 a_1026_45630.t109 7.285
R881 a_1026_45630.n70 a_1026_45630.t177 21.655
R882 a_1026_45630.n69 a_1026_45630.n59 220.884
R883 a_1026_45630.n59 a_1026_45630.n68 7.345
R884 a_1026_45630.n68 a_1026_45630.t89 7.285
R885 a_1026_45630.n68 a_1026_45630.n67 14.37
R886 a_1026_45630.n67 a_1026_45630.t155 7.285
R887 a_1026_45630.n67 a_1026_45630.n66 14.37
R888 a_1026_45630.n66 a_1026_45630.t201 7.285
R889 a_1026_45630.n66 a_1026_45630.n65 14.37
R890 a_1026_45630.n65 a_1026_45630.t67 7.285
R891 a_1026_45630.n65 a_1026_45630.n64 14.395
R892 a_1026_45630.n64 a_1026_45630.t116 7.285
R893 a_1026_45630.n64 a_1026_45630.n63 14.37
R894 a_1026_45630.n63 a_1026_45630.t71 7.285
R895 a_1026_45630.n63 a_1026_45630.n62 14.37
R896 a_1026_45630.n62 a_1026_45630.t139 7.285
R897 a_1026_45630.n62 a_1026_45630.n61 14.37
R898 a_1026_45630.n61 a_1026_45630.t184 7.285
R899 a_1026_45630.n61 a_1026_45630.n60 15.728
R900 a_1026_45630.n60 a_1026_45630.t144 7.285
R901 a_1026_45630.n60 a_1026_45630.t15 21.655
R902 a_1026_45630.n59 a_1026_45630.n49 205.473
R903 a_1026_45630.n49 a_1026_45630.n58 7.345
R904 a_1026_45630.n58 a_1026_45630.t173 7.285
R905 a_1026_45630.n58 a_1026_45630.n57 14.37
R906 a_1026_45630.n57 a_1026_45630.t37 7.285
R907 a_1026_45630.n57 a_1026_45630.n56 14.37
R908 a_1026_45630.n56 a_1026_45630.t87 7.285
R909 a_1026_45630.n56 a_1026_45630.n55 14.37
R910 a_1026_45630.n55 a_1026_45630.t153 7.285
R911 a_1026_45630.n55 a_1026_45630.n54 14.395
R912 a_1026_45630.n54 a_1026_45630.t4 7.285
R913 a_1026_45630.n54 a_1026_45630.n53 14.37
R914 a_1026_45630.n53 a_1026_45630.t157 7.285
R915 a_1026_45630.n53 a_1026_45630.n52 14.37
R916 a_1026_45630.n52 a_1026_45630.t26 7.285
R917 a_1026_45630.n52 a_1026_45630.n51 14.37
R918 a_1026_45630.n51 a_1026_45630.t70 7.285
R919 a_1026_45630.n51 a_1026_45630.n50 15.728
R920 a_1026_45630.n50 a_1026_45630.t182 7.285
R921 a_1026_45630.n50 a_1026_45630.t45 21.655
R922 a_1026_45630.n49 a_1026_45630.n39 228.589
R923 a_1026_45630.n39 a_1026_45630.n48 7.345
R924 a_1026_45630.n48 a_1026_45630.t12 7.285
R925 a_1026_45630.n48 a_1026_45630.n47 14.37
R926 a_1026_45630.n47 a_1026_45630.t77 7.285
R927 a_1026_45630.n47 a_1026_45630.n46 14.37
R928 a_1026_45630.n46 a_1026_45630.t124 7.285
R929 a_1026_45630.n46 a_1026_45630.n45 14.37
R930 a_1026_45630.n45 a_1026_45630.t191 7.285
R931 a_1026_45630.n45 a_1026_45630.n44 14.395
R932 a_1026_45630.n44 a_1026_45630.t43 7.285
R933 a_1026_45630.n44 a_1026_45630.n43 14.37
R934 a_1026_45630.n43 a_1026_45630.t195 7.285
R935 a_1026_45630.n43 a_1026_45630.n42 14.37
R936 a_1026_45630.n42 a_1026_45630.t64 7.285
R937 a_1026_45630.n42 a_1026_45630.n41 14.37
R938 a_1026_45630.n41 a_1026_45630.t112 7.285
R939 a_1026_45630.n41 a_1026_45630.n40 15.728
R940 a_1026_45630.n40 a_1026_45630.t24 7.285
R941 a_1026_45630.n40 a_1026_45630.t95 21.655
R942 a_1026_45630.n39 a_1026_45630.n29 198.41
R943 a_1026_45630.n29 a_1026_45630.n38 7.345
R944 a_1026_45630.n38 a_1026_45630.t49 7.285
R945 a_1026_45630.n38 a_1026_45630.n37 14.37
R946 a_1026_45630.n37 a_1026_45630.t118 7.285
R947 a_1026_45630.n37 a_1026_45630.n36 14.37
R948 a_1026_45630.n36 a_1026_45630.t163 7.285
R949 a_1026_45630.n36 a_1026_45630.n35 14.37
R950 a_1026_45630.n35 a_1026_45630.t30 7.285
R951 a_1026_45630.n35 a_1026_45630.n34 14.395
R952 a_1026_45630.n34 a_1026_45630.t85 7.285
R953 a_1026_45630.n34 a_1026_45630.n33 14.37
R954 a_1026_45630.n33 a_1026_45630.t34 7.285
R955 a_1026_45630.n33 a_1026_45630.n32 14.37
R956 a_1026_45630.n32 a_1026_45630.t107 7.285
R957 a_1026_45630.n32 a_1026_45630.n31 14.37
R958 a_1026_45630.n31 a_1026_45630.t150 7.285
R959 a_1026_45630.n31 a_1026_45630.n30 15.728
R960 a_1026_45630.n30 a_1026_45630.t60 7.285
R961 a_1026_45630.n30 a_1026_45630.t131 21.655
R962 a_1026_45630.n29 a_1026_45630.n20 220.523
R963 a_1026_45630.n28 a_1026_45630.t17 21.655
R964 a_1026_45630.n28 a_1026_45630.t148 7.285
R965 a_1026_45630.n27 a_1026_45630.t33 7.285
R966 a_1026_45630.n27 a_1026_45630.n28 15.728
R967 a_1026_45630.n26 a_1026_45630.t188 7.285
R968 a_1026_45630.n26 a_1026_45630.n27 14.37
R969 a_1026_45630.n25 a_1026_45630.t121 7.285
R970 a_1026_45630.n25 a_1026_45630.n26 14.37
R971 a_1026_45630.n24 a_1026_45630.t170 7.285
R972 a_1026_45630.n24 a_1026_45630.n25 14.37
R973 a_1026_45630.n23 a_1026_45630.t117 7.285
R974 a_1026_45630.n23 a_1026_45630.n24 14.395
R975 a_1026_45630.n22 a_1026_45630.t48 7.285
R976 a_1026_45630.n22 a_1026_45630.n23 14.37
R977 a_1026_45630.n21 a_1026_45630.t5 7.285
R978 a_1026_45630.n21 a_1026_45630.n22 14.37
R979 a_1026_45630.n20 a_1026_45630.t138 7.285
R980 a_1026_45630.n20 a_1026_45630.n21 14.37
R981 a_1026_45630.n119 a_1026_45630.n19 6.95
R982 a_1026_45630.n19 a_1026_45630.t96 7.285
R983 a_1026_45630.n19 a_1026_45630.n18 14.37
R984 a_1026_45630.n18 a_1026_45630.t159 7.285
R985 a_1026_45630.n18 a_1026_45630.n17 14.37
R986 a_1026_45630.n17 a_1026_45630.t6 7.285
R987 a_1026_45630.n17 a_1026_45630.n16 14.37
R988 a_1026_45630.n16 a_1026_45630.t72 7.285
R989 a_1026_45630.n16 a_1026_45630.n15 14.395
R990 a_1026_45630.n15 a_1026_45630.t123 7.285
R991 a_1026_45630.n15 a_1026_45630.n14 14.37
R992 a_1026_45630.n14 a_1026_45630.t76 7.285
R993 a_1026_45630.n14 a_1026_45630.n13 14.37
R994 a_1026_45630.n13 a_1026_45630.t143 7.285
R995 a_1026_45630.n13 a_1026_45630.n12 14.37
R996 a_1026_45630.n12 a_1026_45630.t190 7.285
R997 a_1026_45630.n12 a_1026_45630.n11 15.728
R998 a_1026_45630.n11 a_1026_45630.t105 7.285
R999 a_1026_45630.n11 a_1026_45630.t172 21.655
R1000 a_1026_45630.n200 a_1026_45630.n10 7.345
R1001 a_1026_45630.n10 a_1026_45630.t147 7.285
R1002 a_1026_45630.n10 a_1026_45630.n9 14.37
R1003 a_1026_45630.n9 a_1026_45630.t18 7.285
R1004 a_1026_45630.n9 a_1026_45630.n8 14.37
R1005 a_1026_45630.n8 a_1026_45630.t59 7.285
R1006 a_1026_45630.n8 a_1026_45630.n7 14.37
R1007 a_1026_45630.n7 a_1026_45630.t129 7.285
R1008 a_1026_45630.n7 a_1026_45630.n6 14.395
R1009 a_1026_45630.n6 a_1026_45630.t180 7.285
R1010 a_1026_45630.n6 a_1026_45630.n5 14.37
R1011 a_1026_45630.n5 a_1026_45630.t133 7.285
R1012 a_1026_45630.n5 a_1026_45630.n4 14.37
R1013 a_1026_45630.n4 a_1026_45630.t202 7.285
R1014 a_1026_45630.n4 a_1026_45630.n3 14.37
R1015 a_1026_45630.n3 a_1026_45630.t44 7.285
R1016 a_1026_45630.n3 a_1026_45630.n2 15.728
R1017 a_1026_45630.n2 a_1026_45630.t7 7.285
R1018 a_1026_45630.n2 a_1026_45630.t73 21.655
R1019 Vso1b.t0 Vso1b.n0 17.676
R1020 Vso1b.n0 Vso1b.n3 6.258
R1021 Vso1b.n3 Vso1b.t4 420.019
R1022 Vso1b.n3 Vso1b.n1 157.922
R1023 Vso1b.n1 Vso1b.n2 73.815
R1024 Vso1b.n2 Vso1b.t2 580.661
R1025 Vso1b.n2 Vso1b.t3 185.839
R1026 Vso1b.n1 Vso1b.t5 275.185
R1027 Vso1b.n0 Vso1b.t1 132.095
R1028 a_4226_11420.t0 a_4226_11420.n0 18.871
R1029 a_4226_11420.n0 a_4226_11420.n1 1.803
R1030 a_4226_11420.n1 a_4226_11420.t2 26.764
R1031 a_4226_11420.n1 a_4226_11420.n2 2.933
R1032 a_4226_11420.n2 a_4226_11420.t3 433.701
R1033 a_4226_11420.n2 a_4226_11420.t4 598.416
R1034 a_4226_11420.n0 a_4226_11420.t1 17.028
R1035 a_27962_17218.n4 a_27962_17218.n5 75.708
R1036 a_27962_17218.n0 a_27962_17218.n1 75.707
R1037 a_27962_17218.n1 a_27962_17218.n2 75.707
R1038 a_27962_17218.n2 a_27962_17218.n3 75.707
R1039 a_27962_17218.n3 a_27962_17218.n4 75.707
R1040 a_27962_17218.n6 a_27962_17218.n0 75.707
R1041 a_27962_17218.n4 a_27962_17218.t11 17.401
R1042 a_27962_17218.n3 a_27962_17218.t7 17.401
R1043 a_27962_17218.n2 a_27962_17218.t12 17.401
R1044 a_27962_17218.n1 a_27962_17218.t8 17.401
R1045 a_27962_17218.n0 a_27962_17218.t13 17.401
R1046 a_27962_17218.n5 a_27962_17218.t10 17.4
R1047 a_27962_17218.n5 a_27962_17218.t0 17.4
R1048 a_27962_17218.n4 a_27962_17218.t4 17.4
R1049 a_27962_17218.n3 a_27962_17218.t1 17.4
R1050 a_27962_17218.n2 a_27962_17218.t5 17.4
R1051 a_27962_17218.n1 a_27962_17218.t2 17.4
R1052 a_27962_17218.n0 a_27962_17218.t3 17.4
R1053 a_27962_17218.n6 a_27962_17218.t9 17.4
R1054 a_27962_17218.t6 a_27962_17218.n6 17.4
R1055 a_28220_17218.n0 a_28220_17218.n3 75.439
R1056 a_28220_17218.n4 a_28220_17218.n5 75.437
R1057 a_28220_17218.n2 a_28220_17218.n1 75.436
R1058 a_28220_17218.n3 a_28220_17218.n2 75.436
R1059 a_28220_17218.n1 a_28220_17218.n6 75.436
R1060 a_28220_17218.n0 a_28220_17218.n4 75.435
R1061 a_28220_17218.n0 a_28220_17218.t4 17.401
R1062 a_28220_17218.n4 a_28220_17218.t0 17.401
R1063 a_28220_17218.n3 a_28220_17218.t5 17.401
R1064 a_28220_17218.n2 a_28220_17218.t1 17.401
R1065 a_28220_17218.n1 a_28220_17218.t2 17.401
R1066 a_28220_17218.n5 a_28220_17218.t3 17.4
R1067 a_28220_17218.n5 a_28220_17218.t11 17.4
R1068 a_28220_17218.n4 a_28220_17218.t8 17.4
R1069 a_28220_17218.n3 a_28220_17218.t9 17.4
R1070 a_28220_17218.n2 a_28220_17218.t13 17.4
R1071 a_28220_17218.n1 a_28220_17218.t7 17.4
R1072 a_28220_17218.n6 a_28220_17218.t6 17.4
R1073 a_28220_17218.n6 a_28220_17218.t10 17.4
R1074 a_28220_17218.t12 a_28220_17218.n0 17.4
R1075 a_29252_17218.n4 a_29252_17218.n5 75.708
R1076 a_29252_17218.n0 a_29252_17218.n1 75.707
R1077 a_29252_17218.n1 a_29252_17218.n2 75.707
R1078 a_29252_17218.n2 a_29252_17218.n3 75.707
R1079 a_29252_17218.n3 a_29252_17218.n4 75.707
R1080 a_29252_17218.n6 a_29252_17218.n0 75.707
R1081 a_29252_17218.n4 a_29252_17218.t7 17.401
R1082 a_29252_17218.n3 a_29252_17218.t11 17.401
R1083 a_29252_17218.n2 a_29252_17218.t8 17.401
R1084 a_29252_17218.n1 a_29252_17218.t9 17.401
R1085 a_29252_17218.n0 a_29252_17218.t10 17.401
R1086 a_29252_17218.n5 a_29252_17218.t13 17.4
R1087 a_29252_17218.n5 a_29252_17218.t0 17.4
R1088 a_29252_17218.n4 a_29252_17218.t4 17.4
R1089 a_29252_17218.n3 a_29252_17218.t1 17.4
R1090 a_29252_17218.n2 a_29252_17218.t5 17.4
R1091 a_29252_17218.n1 a_29252_17218.t2 17.4
R1092 a_29252_17218.n0 a_29252_17218.t3 17.4
R1093 a_29252_17218.n6 a_29252_17218.t12 17.4
R1094 a_29252_17218.t6 a_29252_17218.n6 17.4
R1095 a_29510_17218.n0 a_29510_17218.n3 75.71
R1096 a_29510_17218.n4 a_29510_17218.n5 75.708
R1097 a_29510_17218.n2 a_29510_17218.n1 75.707
R1098 a_29510_17218.n3 a_29510_17218.n2 75.707
R1099 a_29510_17218.n1 a_29510_17218.n6 75.707
R1100 a_29510_17218.n0 a_29510_17218.n4 75.706
R1101 a_29510_17218.n0 a_29510_17218.t10 17.401
R1102 a_29510_17218.n4 a_29510_17218.t13 17.401
R1103 a_29510_17218.n3 a_29510_17218.t11 17.401
R1104 a_29510_17218.n2 a_29510_17218.t7 17.401
R1105 a_29510_17218.n1 a_29510_17218.t8 17.401
R1106 a_29510_17218.n5 a_29510_17218.t9 17.4
R1107 a_29510_17218.n5 a_29510_17218.t5 17.4
R1108 a_29510_17218.n4 a_29510_17218.t2 17.4
R1109 a_29510_17218.n3 a_29510_17218.t3 17.4
R1110 a_29510_17218.n2 a_29510_17218.t0 17.4
R1111 a_29510_17218.n1 a_29510_17218.t1 17.4
R1112 a_29510_17218.n6 a_29510_17218.t12 17.4
R1113 a_29510_17218.n6 a_29510_17218.t4 17.4
R1114 a_29510_17218.t6 a_29510_17218.n0 17.4
R1115 Fvco_By4_QPH.t10 Fvco_By4_QPH.t19 731.89
R1116 Fvco_By4_QPH.t14 Fvco_By4_QPH.t6 731.89
R1117 Fvco_By4_QPH.t3 Fvco_By4_QPH.t13 731.89
R1118 Fvco_By4_QPH.t5 Fvco_By4_QPH.t16 718.506
R1119 Fvco_By4_QPH.t11 Fvco_By4_QPH.t15 710.965
R1120 Fvco_By4_QPH.t7 Fvco_By4_QPH.t14 622.637
R1121 Fvco_By4_QPH.n7 Fvco_By4_QPH.n6 617.524
R1122 Fvco_By4_QPH.n3 Fvco_By4_QPH.n2 580.872
R1123 Fvco_By4_QPH.t15 Fvco_By4_QPH.t2 579.889
R1124 Fvco_By4_QPH.n2 Fvco_By4_QPH.t12 491.229
R1125 Fvco_By4_QPH.n3 Fvco_By4_QPH.t4 489.182
R1126 Fvco_By4_QPH.n8 Fvco_By4_QPH.t11 418.965
R1127 Fvco_By4_QPH.n7 Fvco_By4_QPH.t18 414.13
R1128 Fvco_By4_QPH.n4 Fvco_By4_QPH.t9 349.273
R1129 Fvco_By4_QPH.n1 Fvco_By4_QPH.t8 333.651
R1130 Fvco_By4_QPH.n5 Fvco_By4_QPH.t3 317.894
R1131 Fvco_By4_QPH.n1 Fvco_By4_QPH.t17 297.233
R1132 Fvco_By4_QPH.n5 Fvco_By4_QPH.t5 291.323
R1133 Fvco_By4_QPH.n4 Fvco_By4_QPH.t10 252.624
R1134 Fvco_By4_QPH.n2 Fvco_By4_QPH.t7 227.612
R1135 Fvco_By4_QPH.t9 Fvco_By4_QPH.n3 227.612
R1136 Fvco_By4_QPH.n6 Fvco_By4_QPH.n4 198.896
R1137 Fvco_By4_QPH.n8 Fvco_By4_QPH.n7 152.778
R1138 Fvco_By4_QPH.n0 Fvco_By4_QPH.t0 92.046
R1139 Fvco_By4_QPH.n0 Fvco_By4_QPH.n1 70.221
R1140 Fvco_By4_QPH.n0 Fvco_By4_QPH.t1 61.427
R1141 Fvco_By4_QPH Fvco_By4_QPH.n8 38.508
R1142 Fvco_By4_QPH.n6 Fvco_By4_QPH.n5 31.687
R1143 Fvco_By4_QPH Fvco_By4_QPH.n0 11.126
R1144 a_55602_11692.t0 a_55602_11692.n0 14.504
R1145 a_55602_11692.n0 a_55602_11692.n1 0.395
R1146 a_55602_11692.n0 a_55602_11692.n3 815.609
R1147 a_55602_11692.n3 a_55602_11692.n9 328.781
R1148 a_55602_11692.n10 a_55602_11692.t8 212.622
R1149 a_55602_11692.n11 a_55602_11692.n10 208.271
R1150 a_55602_11692.n9 a_55602_11692.n11 76.046
R1151 a_55602_11692.n11 a_55602_11692.t10 4.351
R1152 a_55602_11692.n10 a_55602_11692.t2 4.351
R1153 a_55602_11692.n5 a_55602_11692.n6 0.001
R1154 a_55602_11692.n7 a_55602_11692.n8 0.001
R1155 a_55602_11692.n5 a_55602_11692.n4 208.271
R1156 a_55602_11692.n7 a_55602_11692.n5 208.271
R1157 a_55602_11692.n9 a_55602_11692.n7 155.811
R1158 a_55602_11692.n8 a_55602_11692.t12 4.35
R1159 a_55602_11692.n8 a_55602_11692.t11 4.35
R1160 a_55602_11692.n6 a_55602_11692.t9 4.35
R1161 a_55602_11692.n6 a_55602_11692.t7 4.35
R1162 a_55602_11692.n4 a_55602_11692.t4 4.35
R1163 a_55602_11692.n4 a_55602_11692.t3 4.35
R1164 a_55602_11692.n3 a_55602_11692.t13 5.714
R1165 a_55602_11692.n1 a_55602_11692.n2 2.815
R1166 a_55602_11692.n2 a_55602_11692.t5 17.453
R1167 a_55602_11692.n2 a_55602_11692.t1 17.451
R1168 a_55602_11692.n1 a_55602_11692.t6 14.331
R1169 a_50320_14126.t0 a_50320_14126.n0 14.302
R1170 a_50320_14126.n7 a_50320_14126.t1 18.036
R1171 a_50320_14126.n0 a_50320_14126.n7 1.885
R1172 a_50320_14126.n7 a_50320_14126.t2 17.538
R1173 a_50320_14126.n0 a_50320_14126.n6 3.212
R1174 a_50320_14126.n6 a_50320_14126.t3 15.994
R1175 a_50320_14126.n6 a_50320_14126.n4 425.295
R1176 a_50320_14126.n5 a_50320_14126.t9 48.21
R1177 a_50320_14126.n5 a_50320_14126.t4 127.084
R1178 a_50320_14126.n4 a_50320_14126.n5 1.418
R1179 a_50320_14126.n4 a_50320_14126.n2 31.793
R1180 a_50320_14126.n3 a_50320_14126.t6 48.21
R1181 a_50320_14126.n3 a_50320_14126.t8 127.084
R1182 a_50320_14126.n2 a_50320_14126.n3 1.418
R1183 a_50320_14126.n1 a_50320_14126.t5 48.21
R1184 a_50320_14126.n1 a_50320_14126.t7 127.084
R1185 a_50320_14126.n2 a_50320_14126.n1 35.06
R1186 a_49874_4150.t1 a_49874_4150.t0 40.008
R1187 a_54950_4814.t0 a_54950_4814.t1 27.186
R1188 a_14188_14050.t12 a_14188_14050.t52 1273.78
R1189 a_14188_14050.t12 a_14188_14050.t31 161.992
R1190 a_14188_14050.t31 a_14188_14050.t39 126.193
R1191 a_14188_14050.t31 a_14188_14050.t49 113.753
R1192 a_14188_14050.t31 a_14188_14050.t46 113.753
R1193 a_14188_14050.t31 a_14188_14050.t11 113.753
R1194 a_14188_14050.t31 a_14188_14050.t23 113.753
R1195 a_14188_14050.t31 a_14188_14050.t6 113.753
R1196 a_14188_14050.t31 a_14188_14050.t18 113.753
R1197 a_14188_14050.t31 a_14188_14050.t40 113.753
R1198 a_14188_14050.t31 a_14188_14050.t54 113.753
R1199 a_14188_14050.t31 a_14188_14050.t9 113.753
R1200 a_14188_14050.t31 a_14188_14050.t8 113.753
R1201 a_14188_14050.t31 a_14188_14050.t26 113.753
R1202 a_14188_14050.t31 a_14188_14050.t41 113.753
R1203 a_14188_14050.t31 a_14188_14050.t24 113.753
R1204 a_14188_14050.t31 a_14188_14050.t38 113.753
R1205 a_14188_14050.t31 a_14188_14050.t56 113.753
R1206 a_14188_14050.t31 a_14188_14050.t21 113.753
R1207 a_14188_14050.t31 a_14188_14050.t36 113.753
R1208 a_14188_14050.t31 a_14188_14050.t33 113.753
R1209 a_14188_14050.t31 a_14188_14050.t55 113.753
R1210 a_14188_14050.t31 a_14188_14050.t10 113.753
R1211 a_14188_14050.t31 a_14188_14050.t50 113.753
R1212 a_14188_14050.t31 a_14188_14050.t5 113.753
R1213 a_14188_14050.t31 a_14188_14050.t25 113.753
R1214 a_14188_14050.t31 a_14188_14050.t48 113.753
R1215 a_14188_14050.t31 a_14188_14050.t4 113.753
R1216 a_14188_14050.t31 a_14188_14050.t59 113.753
R1217 a_14188_14050.t31 a_14188_14050.t22 113.753
R1218 a_14188_14050.t31 a_14188_14050.t37 113.753
R1219 a_14188_14050.t31 a_14188_14050.t19 113.753
R1220 a_14188_14050.t31 a_14188_14050.t30 113.753
R1221 a_14188_14050.t31 a_14188_14050.t53 113.753
R1222 a_14188_14050.t31 a_14188_14050.t2 113.753
R1223 a_14188_14050.t31 a_14188_14050.t15 113.753
R1224 a_14188_14050.t31 a_14188_14050.t14 113.753
R1225 a_14188_14050.t31 a_14188_14050.t35 113.753
R1226 a_14188_14050.t31 a_14188_14050.t47 113.753
R1227 a_14188_14050.t31 a_14188_14050.t29 113.753
R1228 a_14188_14050.t31 a_14188_14050.t44 113.753
R1229 a_14188_14050.t31 a_14188_14050.t7 113.753
R1230 a_14188_14050.t31 a_14188_14050.t45 113.753
R1231 a_14188_14050.t31 a_14188_14050.t60 113.753
R1232 a_14188_14050.t31 a_14188_14050.t58 113.753
R1233 a_14188_14050.t31 a_14188_14050.t20 113.753
R1234 a_14188_14050.t31 a_14188_14050.t28 113.753
R1235 a_14188_14050.t31 a_14188_14050.t43 113.753
R1236 a_14188_14050.t31 a_14188_14050.t42 113.753
R1237 a_14188_14050.t31 a_14188_14050.t3 113.753
R1238 a_14188_14050.t31 a_14188_14050.t16 113.753
R1239 a_14188_14050.t31 a_14188_14050.t57 113.753
R1240 a_14188_14050.t31 a_14188_14050.t13 113.753
R1241 a_14188_14050.t31 a_14188_14050.t32 113.753
R1242 a_14188_14050.t31 a_14188_14050.t34 113.753
R1243 a_14188_14050.t31 a_14188_14050.t17 113.753
R1244 a_14188_14050.t31 a_14188_14050.t27 113.753
R1245 a_14188_14050.t31 a_14188_14050.t51 113.753
R1246 a_14188_14050.t12 a_14188_14050.t0 57.908
R1247 a_14188_14050.t1 a_14188_14050.t12 57.821
R1248 a_22629_5596.n0 a_22629_5596.n1 75.71
R1249 a_22629_5596.n4 a_22629_5596.n5 75.708
R1250 a_22629_5596.n2 a_22629_5596.n3 75.707
R1251 a_22629_5596.n3 a_22629_5596.n4 75.707
R1252 a_22629_5596.n1 a_22629_5596.n6 75.707
R1253 a_22629_5596.n0 a_22629_5596.n2 75.706
R1254 a_22629_5596.n0 a_22629_5596.t10 17.401
R1255 a_22629_5596.n4 a_22629_5596.t11 17.401
R1256 a_22629_5596.n3 a_22629_5596.t13 17.401
R1257 a_22629_5596.n2 a_22629_5596.t9 17.401
R1258 a_22629_5596.n1 a_22629_5596.t12 17.401
R1259 a_22629_5596.n5 a_22629_5596.t8 17.4
R1260 a_22629_5596.n5 a_22629_5596.t3 17.4
R1261 a_22629_5596.n4 a_22629_5596.t0 17.4
R1262 a_22629_5596.n3 a_22629_5596.t5 17.4
R1263 a_22629_5596.n2 a_22629_5596.t1 17.4
R1264 a_22629_5596.n1 a_22629_5596.t4 17.4
R1265 a_22629_5596.n6 a_22629_5596.t7 17.4
R1266 a_22629_5596.n6 a_22629_5596.t2 17.4
R1267 a_22629_5596.t6 a_22629_5596.n0 17.4
R1268 a_23145_5596.n0 a_23145_5596.n2 75.71
R1269 a_23145_5596.n4 a_23145_5596.n5 75.708
R1270 a_23145_5596.n2 a_23145_5596.n1 75.707
R1271 a_23145_5596.n3 a_23145_5596.n4 75.707
R1272 a_23145_5596.n1 a_23145_5596.n6 75.707
R1273 a_23145_5596.n0 a_23145_5596.n3 75.706
R1274 a_23145_5596.n0 a_23145_5596.t7 17.401
R1275 a_23145_5596.n4 a_23145_5596.t6 17.401
R1276 a_23145_5596.n3 a_23145_5596.t4 17.401
R1277 a_23145_5596.n2 a_23145_5596.t5 17.401
R1278 a_23145_5596.n1 a_23145_5596.t1 17.401
R1279 a_23145_5596.n5 a_23145_5596.t3 17.4
R1280 a_23145_5596.n5 a_23145_5596.t13 17.4
R1281 a_23145_5596.n4 a_23145_5596.t11 17.4
R1282 a_23145_5596.n3 a_23145_5596.t9 17.4
R1283 a_23145_5596.n2 a_23145_5596.t10 17.4
R1284 a_23145_5596.n1 a_23145_5596.t8 17.4
R1285 a_23145_5596.n6 a_23145_5596.t2 17.4
R1286 a_23145_5596.n6 a_23145_5596.t12 17.4
R1287 a_23145_5596.t0 a_23145_5596.n0 17.4
R1288 a_23403_5596.n6 a_23403_5596.n4 75.711
R1289 a_23403_5596.n1 a_23403_5596.n0 75.707
R1290 a_23403_5596.n2 a_23403_5596.n1 75.707
R1291 a_23403_5596.n3 a_23403_5596.n2 75.707
R1292 a_23403_5596.n4 a_23403_5596.n3 75.707
R1293 a_23403_5596.n0 a_23403_5596.n5 75.707
R1294 a_23403_5596.n4 a_23403_5596.t6 17.401
R1295 a_23403_5596.n3 a_23403_5596.t4 17.401
R1296 a_23403_5596.n2 a_23403_5596.t2 17.401
R1297 a_23403_5596.n1 a_23403_5596.t5 17.401
R1298 a_23403_5596.n0 a_23403_5596.t1 17.401
R1299 a_23403_5596.n4 a_23403_5596.t9 17.4
R1300 a_23403_5596.n3 a_23403_5596.t7 17.4
R1301 a_23403_5596.n2 a_23403_5596.t10 17.4
R1302 a_23403_5596.n1 a_23403_5596.t8 17.4
R1303 a_23403_5596.n0 a_23403_5596.t13 17.4
R1304 a_23403_5596.n5 a_23403_5596.t3 17.4
R1305 a_23403_5596.n5 a_23403_5596.t11 17.4
R1306 a_23403_5596.n6 a_23403_5596.t0 17.4
R1307 a_23403_5596.t12 a_23403_5596.n6 17.4
R1308 a_53292_4814.t0 a_53292_4814.t1 27.186
R1309 a_22887_5596.n0 a_22887_5596.n2 75.439
R1310 a_22887_5596.n4 a_22887_5596.n5 75.437
R1311 a_22887_5596.n2 a_22887_5596.n1 75.436
R1312 a_22887_5596.n3 a_22887_5596.n4 75.436
R1313 a_22887_5596.n1 a_22887_5596.n6 75.436
R1314 a_22887_5596.n0 a_22887_5596.n3 75.435
R1315 a_22887_5596.n0 a_22887_5596.t7 17.401
R1316 a_22887_5596.n4 a_22887_5596.t13 17.401
R1317 a_22887_5596.n3 a_22887_5596.t11 17.401
R1318 a_22887_5596.n2 a_22887_5596.t12 17.401
R1319 a_22887_5596.n1 a_22887_5596.t10 17.401
R1320 a_22887_5596.n5 a_22887_5596.t9 17.4
R1321 a_22887_5596.n5 a_22887_5596.t1 17.4
R1322 a_22887_5596.n4 a_22887_5596.t5 17.4
R1323 a_22887_5596.n3 a_22887_5596.t3 17.4
R1324 a_22887_5596.n2 a_22887_5596.t4 17.4
R1325 a_22887_5596.n1 a_22887_5596.t2 17.4
R1326 a_22887_5596.n6 a_22887_5596.t8 17.4
R1327 a_22887_5596.n6 a_22887_5596.t0 17.4
R1328 a_22887_5596.t6 a_22887_5596.n0 17.4
R1329 a_26036_4988.t16 a_26036_4988.t22 1273.78
R1330 a_26036_4988.t16 a_26036_4988.t20 415.476
R1331 a_26036_4988.t20 a_26036_4988.t8 127.909
R1332 a_26036_4988.t20 a_26036_4988.t37 113.753
R1333 a_26036_4988.t20 a_26036_4988.t34 113.753
R1334 a_26036_4988.t20 a_26036_4988.t32 113.753
R1335 a_26036_4988.t20 a_26036_4988.t45 113.753
R1336 a_26036_4988.t20 a_26036_4988.t7 113.753
R1337 a_26036_4988.t20 a_26036_4988.t4 113.753
R1338 a_26036_4988.t20 a_26036_4988.t60 113.753
R1339 a_26036_4988.t20 a_26036_4988.t14 113.753
R1340 a_26036_4988.t20 a_26036_4988.t46 113.753
R1341 a_26036_4988.t20 a_26036_4988.t10 113.753
R1342 a_26036_4988.t20 a_26036_4988.t6 113.753
R1343 a_26036_4988.t20 a_26036_4988.t3 113.753
R1344 a_26036_4988.t20 a_26036_4988.t15 113.753
R1345 a_26036_4988.t20 a_26036_4988.t41 113.753
R1346 a_26036_4988.t20 a_26036_4988.t38 113.753
R1347 a_26036_4988.t20 a_26036_4988.t35 113.753
R1348 a_26036_4988.t20 a_26036_4988.t54 113.753
R1349 a_26036_4988.t20 a_26036_4988.t51 113.753
R1350 a_26036_4988.t20 a_26036_4988.t48 113.753
R1351 a_26036_4988.t20 a_26036_4988.t5 113.753
R1352 a_26036_4988.t20 a_26036_4988.t27 113.753
R1353 a_26036_4988.t20 a_26036_4988.t24 113.753
R1354 a_26036_4988.t20 a_26036_4988.t18 113.753
R1355 a_26036_4988.t20 a_26036_4988.t36 113.753
R1356 a_26036_4988.t20 a_26036_4988.t29 113.753
R1357 a_26036_4988.t20 a_26036_4988.t26 113.753
R1358 a_26036_4988.t20 a_26036_4988.t23 113.753
R1359 a_26036_4988.t20 a_26036_4988.t39 113.753
R1360 a_26036_4988.t20 a_26036_4988.t58 113.753
R1361 a_26036_4988.t20 a_26036_4988.t56 113.753
R1362 a_26036_4988.t20 a_26036_4988.t52 113.753
R1363 a_26036_4988.t20 a_26036_4988.t59 113.753
R1364 a_26036_4988.t20 a_26036_4988.t57 113.753
R1365 a_26036_4988.t20 a_26036_4988.t55 113.753
R1366 a_26036_4988.t20 a_26036_4988.t11 113.753
R1367 a_26036_4988.t20 a_26036_4988.t31 113.753
R1368 a_26036_4988.t20 a_26036_4988.t30 113.753
R1369 a_26036_4988.t20 a_26036_4988.t28 113.753
R1370 a_26036_4988.t20 a_26036_4988.t42 113.753
R1371 a_26036_4988.t20 a_26036_4988.t19 113.753
R1372 a_26036_4988.t20 a_26036_4988.t44 113.753
R1373 a_26036_4988.t20 a_26036_4988.t43 113.753
R1374 a_26036_4988.t20 a_26036_4988.t40 113.753
R1375 a_26036_4988.t20 a_26036_4988.t49 113.753
R1376 a_26036_4988.t20 a_26036_4988.t13 113.753
R1377 a_26036_4988.t20 a_26036_4988.t12 113.753
R1378 a_26036_4988.t20 a_26036_4988.t9 113.753
R1379 a_26036_4988.t20 a_26036_4988.t33 113.753
R1380 a_26036_4988.t20 a_26036_4988.t53 113.753
R1381 a_26036_4988.t20 a_26036_4988.t50 113.753
R1382 a_26036_4988.t20 a_26036_4988.t47 113.753
R1383 a_26036_4988.t20 a_26036_4988.t2 113.753
R1384 a_26036_4988.t20 a_26036_4988.t25 113.753
R1385 a_26036_4988.t20 a_26036_4988.t21 113.753
R1386 a_26036_4988.t20 a_26036_4988.t17 113.753
R1387 a_26036_4988.t0 a_26036_4988.t16 81.094
R1388 a_26036_4988.t16 a_26036_4988.t1 33.947
R1389 a_28736_5597.n4 a_28736_5597.n5 75.708
R1390 a_28736_5597.n0 a_28736_5597.n1 75.707
R1391 a_28736_5597.n1 a_28736_5597.n2 75.707
R1392 a_28736_5597.n2 a_28736_5597.n3 75.707
R1393 a_28736_5597.n3 a_28736_5597.n4 75.707
R1394 a_28736_5597.n6 a_28736_5597.n0 75.707
R1395 a_28736_5597.n4 a_28736_5597.t3 17.401
R1396 a_28736_5597.n3 a_28736_5597.t12 17.401
R1397 a_28736_5597.n2 a_28736_5597.t9 17.401
R1398 a_28736_5597.n1 a_28736_5597.t2 17.401
R1399 a_28736_5597.n0 a_28736_5597.t11 17.401
R1400 a_28736_5597.n5 a_28736_5597.t13 17.4
R1401 a_28736_5597.n5 a_28736_5597.t1 17.4
R1402 a_28736_5597.n4 a_28736_5597.t4 17.4
R1403 a_28736_5597.n3 a_28736_5597.t7 17.4
R1404 a_28736_5597.n2 a_28736_5597.t5 17.4
R1405 a_28736_5597.n1 a_28736_5597.t8 17.4
R1406 a_28736_5597.n0 a_28736_5597.t6 17.4
R1407 a_28736_5597.n6 a_28736_5597.t10 17.4
R1408 a_28736_5597.t0 a_28736_5597.n6 17.4
R1409 a_28994_5597.n4 a_28994_5597.n5 75.708
R1410 a_28994_5597.n0 a_28994_5597.n1 75.707
R1411 a_28994_5597.n1 a_28994_5597.n2 75.707
R1412 a_28994_5597.n2 a_28994_5597.n3 75.707
R1413 a_28994_5597.n3 a_28994_5597.n4 75.707
R1414 a_28994_5597.n6 a_28994_5597.n0 75.707
R1415 a_28994_5597.n4 a_28994_5597.t8 17.401
R1416 a_28994_5597.n3 a_28994_5597.t11 17.401
R1417 a_28994_5597.n2 a_28994_5597.t9 17.401
R1418 a_28994_5597.n1 a_28994_5597.t7 17.401
R1419 a_28994_5597.n0 a_28994_5597.t13 17.401
R1420 a_28994_5597.n5 a_28994_5597.t12 17.4
R1421 a_28994_5597.n5 a_28994_5597.t0 17.4
R1422 a_28994_5597.n4 a_28994_5597.t4 17.4
R1423 a_28994_5597.n3 a_28994_5597.t2 17.4
R1424 a_28994_5597.n2 a_28994_5597.t5 17.4
R1425 a_28994_5597.n1 a_28994_5597.t3 17.4
R1426 a_28994_5597.n0 a_28994_5597.t1 17.4
R1427 a_28994_5597.n6 a_28994_5597.t10 17.4
R1428 a_28994_5597.t6 a_28994_5597.n6 17.4
R1429 CLK_BY_4_IPH.n0 CLK_BY_4_IPH.t4 440.519
R1430 CLK_BY_4_IPH.n0 CLK_BY_4_IPH.t3 402.739
R1431 CLK_BY_4_IPH.n2 CLK_BY_4_IPH.t2 227.612
R1432 CLK_BY_4_IPH.n1 CLK_BY_4_IPH.t1 227.612
R1433 CLK_BY_4_IPH.n3 CLK_BY_4_IPH.n2 195.608
R1434 CLK_BY_4_IPH.n1 CLK_BY_4_IPH.n0 183.872
R1435 CLK_BY_4_IPH.n2 CLK_BY_4_IPH.n1 45.046
R1436 CLK_BY_4_IPH.n3 CLK_BY_4_IPH.t0 40.317
R1437 CLK_BY_4_IPH CLK_BY_4_IPH.n3 11.83
R1438 vctrl.t0 vctrl.n0 16.252
R1439 vctrl.n0 vctrl.t2 16.252
R1440 vctrl.n2 vctrl.n1 0.275
R1441 vctrl.n1 vctrl.n0 2.303
R1442 vctrl.n1 vctrl.t1 24.647
R1443 vctrl vctrl.n2 41.937
R1444 vctrl vctrl.n3 1.429
R1445 vctrl.n3 vctrl.n4 0.561
R1446 vctrl.n4 vctrl.t6 0.589
R1447 vctrl.n4 vctrl.t5 0.028
R1448 vctrl.n3 vctrl.t4 0.028
R1449 vctrl.n2 vctrl.t3 24.662
R1450 a_25099_11445.t52 a_25099_11445.t40 1273.78
R1451 a_25099_11445.t52 a_25099_11445.t15 218.051
R1452 a_25099_11445.t15 a_25099_11445.t20 127.858
R1453 a_25099_11445.t15 a_25099_11445.t48 113.753
R1454 a_25099_11445.t15 a_25099_11445.t8 113.753
R1455 a_25099_11445.t15 a_25099_11445.t29 113.753
R1456 a_25099_11445.t15 a_25099_11445.t21 113.753
R1457 a_25099_11445.t15 a_25099_11445.t41 113.753
R1458 a_25099_11445.t15 a_25099_11445.t58 113.753
R1459 a_25099_11445.t15 a_25099_11445.t56 113.753
R1460 a_25099_11445.t15 a_25099_11445.t6 113.753
R1461 a_25099_11445.t15 a_25099_11445.t16 113.753
R1462 a_25099_11445.t15 a_25099_11445.t37 113.753
R1463 a_25099_11445.t15 a_25099_11445.t53 113.753
R1464 a_25099_11445.t15 a_25099_11445.t19 113.753
R1465 a_25099_11445.t15 a_25099_11445.t50 113.753
R1466 a_25099_11445.t15 a_25099_11445.t10 113.753
R1467 a_25099_11445.t15 a_25099_11445.t31 113.753
R1468 a_25099_11445.t15 a_25099_11445.t26 113.753
R1469 a_25099_11445.t15 a_25099_11445.t35 113.753
R1470 a_25099_11445.t15 a_25099_11445.t46 113.753
R1471 a_25099_11445.t15 a_25099_11445.t4 113.753
R1472 a_25099_11445.t15 a_25099_11445.t23 113.753
R1473 a_25099_11445.t15 a_25099_11445.t42 113.753
R1474 a_25099_11445.t15 a_25099_11445.t59 113.753
R1475 a_25099_11445.t15 a_25099_11445.t57 113.753
R1476 a_25099_11445.t15 a_25099_11445.t7 113.753
R1477 a_25099_11445.t15 a_25099_11445.t17 113.753
R1478 a_25099_11445.t15 a_25099_11445.t38 113.753
R1479 a_25099_11445.t15 a_25099_11445.t54 113.753
R1480 a_25099_11445.t15 a_25099_11445.t51 113.753
R1481 a_25099_11445.t15 a_25099_11445.t11 113.753
R1482 a_25099_11445.t15 a_25099_11445.t32 113.753
R1483 a_25099_11445.t15 a_25099_11445.t27 113.753
R1484 a_25099_11445.t15 a_25099_11445.t36 113.753
R1485 a_25099_11445.t15 a_25099_11445.t47 113.753
R1486 a_25099_11445.t15 a_25099_11445.t5 113.753
R1487 a_25099_11445.t15 a_25099_11445.t24 113.753
R1488 a_25099_11445.t15 a_25099_11445.t39 113.753
R1489 a_25099_11445.t15 a_25099_11445.t55 113.753
R1490 a_25099_11445.t15 a_25099_11445.t12 113.753
R1491 a_25099_11445.t15 a_25099_11445.t43 113.753
R1492 a_25099_11445.t15 a_25099_11445.t60 113.753
R1493 a_25099_11445.t15 a_25099_11445.t14 113.753
R1494 a_25099_11445.t15 a_25099_11445.t13 113.753
R1495 a_25099_11445.t15 a_25099_11445.t28 113.753
R1496 a_25099_11445.t15 a_25099_11445.t49 113.753
R1497 a_25099_11445.t15 a_25099_11445.t9 113.753
R1498 a_25099_11445.t15 a_25099_11445.t30 113.753
R1499 a_25099_11445.t15 a_25099_11445.t25 113.753
R1500 a_25099_11445.t15 a_25099_11445.t34 113.753
R1501 a_25099_11445.t15 a_25099_11445.t45 113.753
R1502 a_25099_11445.t15 a_25099_11445.t3 113.753
R1503 a_25099_11445.t15 a_25099_11445.t22 113.753
R1504 a_25099_11445.t15 a_25099_11445.t33 113.753
R1505 a_25099_11445.t15 a_25099_11445.t44 113.753
R1506 a_25099_11445.t15 a_25099_11445.t2 113.753
R1507 a_25099_11445.t15 a_25099_11445.t18 113.753
R1508 a_25099_11445.t1 a_25099_11445.t52 56.779
R1509 a_25099_11445.t52 a_25099_11445.t0 37.09
R1510 a_26589_11500.n0 a_26589_11500.n6 75.709
R1511 a_26589_11500.n4 a_26589_11500.n5 75.708
R1512 a_26589_11500.n1 a_26589_11500.n2 75.707
R1513 a_26589_11500.n2 a_26589_11500.n3 75.707
R1514 a_26589_11500.n3 a_26589_11500.n4 75.707
R1515 a_26589_11500.n0 a_26589_11500.n1 75.706
R1516 a_26589_11500.n0 a_26589_11500.t9 17.401
R1517 a_26589_11500.n4 a_26589_11500.t11 17.401
R1518 a_26589_11500.n3 a_26589_11500.t13 17.401
R1519 a_26589_11500.n2 a_26589_11500.t8 17.401
R1520 a_26589_11500.n1 a_26589_11500.t10 17.401
R1521 a_26589_11500.n5 a_26589_11500.t12 17.4
R1522 a_26589_11500.n5 a_26589_11500.t4 17.4
R1523 a_26589_11500.n4 a_26589_11500.t2 17.4
R1524 a_26589_11500.n3 a_26589_11500.t5 17.4
R1525 a_26589_11500.n2 a_26589_11500.t3 17.4
R1526 a_26589_11500.n1 a_26589_11500.t6 17.4
R1527 a_26589_11500.n6 a_26589_11500.t7 17.4
R1528 a_26589_11500.n6 a_26589_11500.t1 17.4
R1529 a_26589_11500.t0 a_26589_11500.n0 17.4
R1530 a_26847_11500.n4 a_26847_11500.n5 75.708
R1531 a_26847_11500.n0 a_26847_11500.n1 75.707
R1532 a_26847_11500.n1 a_26847_11500.n2 75.707
R1533 a_26847_11500.n2 a_26847_11500.n3 75.707
R1534 a_26847_11500.n3 a_26847_11500.n4 75.707
R1535 a_26847_11500.n6 a_26847_11500.n0 75.707
R1536 a_26847_11500.n4 a_26847_11500.t8 17.401
R1537 a_26847_11500.n3 a_26847_11500.t9 17.401
R1538 a_26847_11500.n2 a_26847_11500.t12 17.401
R1539 a_26847_11500.n1 a_26847_11500.t7 17.401
R1540 a_26847_11500.n0 a_26847_11500.t13 17.401
R1541 a_26847_11500.n5 a_26847_11500.t11 17.4
R1542 a_26847_11500.n5 a_26847_11500.t0 17.4
R1543 a_26847_11500.n4 a_26847_11500.t3 17.4
R1544 a_26847_11500.n3 a_26847_11500.t1 17.4
R1545 a_26847_11500.n2 a_26847_11500.t4 17.4
R1546 a_26847_11500.n1 a_26847_11500.t2 17.4
R1547 a_26847_11500.n0 a_26847_11500.t5 17.4
R1548 a_26847_11500.n6 a_26847_11500.t10 17.4
R1549 a_26847_11500.t6 a_26847_11500.n6 17.4
R1550 a_66154_26414.t0 a_66154_26414.t1 126.642
R1551 a_23919_5596.n0 a_23919_5596.n3 75.71
R1552 a_23919_5596.n4 a_23919_5596.n5 75.708
R1553 a_23919_5596.n2 a_23919_5596.n1 75.707
R1554 a_23919_5596.n3 a_23919_5596.n2 75.707
R1555 a_23919_5596.n1 a_23919_5596.n6 75.707
R1556 a_23919_5596.n0 a_23919_5596.n4 75.706
R1557 a_23919_5596.n0 a_23919_5596.t8 17.401
R1558 a_23919_5596.n4 a_23919_5596.t12 17.401
R1559 a_23919_5596.n3 a_23919_5596.t13 17.401
R1560 a_23919_5596.n2 a_23919_5596.t9 17.401
R1561 a_23919_5596.n1 a_23919_5596.t7 17.401
R1562 a_23919_5596.n5 a_23919_5596.t11 17.4
R1563 a_23919_5596.n5 a_23919_5596.t4 17.4
R1564 a_23919_5596.n4 a_23919_5596.t5 17.4
R1565 a_23919_5596.n3 a_23919_5596.t6 17.4
R1566 a_23919_5596.n2 a_23919_5596.t1 17.4
R1567 a_23919_5596.n1 a_23919_5596.t2 17.4
R1568 a_23919_5596.n6 a_23919_5596.t10 17.4
R1569 a_23919_5596.n6 a_23919_5596.t3 17.4
R1570 a_23919_5596.t0 a_23919_5596.n0 17.4
R1571 a_24177_5596.n0 a_24177_5596.n3 75.71
R1572 a_24177_5596.n4 a_24177_5596.n5 75.708
R1573 a_24177_5596.n2 a_24177_5596.n1 75.707
R1574 a_24177_5596.n3 a_24177_5596.n2 75.707
R1575 a_24177_5596.n1 a_24177_5596.n6 75.707
R1576 a_24177_5596.n0 a_24177_5596.n4 75.706
R1577 a_24177_5596.n0 a_24177_5596.t2 17.401
R1578 a_24177_5596.n4 a_24177_5596.t13 17.401
R1579 a_24177_5596.n3 a_24177_5596.t0 17.401
R1580 a_24177_5596.n2 a_24177_5596.t3 17.401
R1581 a_24177_5596.n1 a_24177_5596.t5 17.401
R1582 a_24177_5596.n5 a_24177_5596.t4 17.4
R1583 a_24177_5596.n5 a_24177_5596.t10 17.4
R1584 a_24177_5596.n4 a_24177_5596.t7 17.4
R1585 a_24177_5596.n3 a_24177_5596.t8 17.4
R1586 a_24177_5596.n2 a_24177_5596.t6 17.4
R1587 a_24177_5596.n1 a_24177_5596.t11 17.4
R1588 a_24177_5596.n6 a_24177_5596.t1 17.4
R1589 a_24177_5596.n6 a_24177_5596.t9 17.4
R1590 a_24177_5596.t12 a_24177_5596.n0 17.4
R1591 a_17685_3840.n29 a_17685_3840.n28 660.793
R1592 a_17685_3840.n57 a_17685_3840.n56 649.743
R1593 a_17685_3840.n60 a_17685_3840.n59 574.593
R1594 a_17685_3840.n30 a_17685_3840.n29 416.406
R1595 a_17685_3840.n61 a_17685_3840.n60 415.789
R1596 a_17685_3840.n26 a_17685_3840.n25 270.636
R1597 a_17685_3840.n28 a_17685_3840.n27 262.3
R1598 a_17685_3840.n29 a_17685_3840.n26 198.935
R1599 a_17685_3840.n59 a_17685_3840.t3 197.212
R1600 a_17685_3840.n27 a_17685_3840.t12 185.816
R1601 a_17685_3840.n28 a_17685_3840.t2 176.327
R1602 a_17685_3840.n58 a_17685_3840.t1 173.989
R1603 a_17685_3840.n26 a_17685_3840.t6 154.605
R1604 a_17685_3840.n25 a_17685_3840.t0 151.674
R1605 a_17685_3840.n62 a_17685_3840.t5 118.032
R1606 a_17685_3840.n60 a_17685_3840.n58 107.97
R1607 a_17685_3840.n31 a_17685_3840.n30 104.297
R1608 a_17685_3840.n63 a_17685_3840.n62 103.649
R1609 a_17685_3840.n67 a_17685_3840.n66 100.879
R1610 a_17685_3840.n64 a_17685_3840.n63 83.404
R1611 a_17685_3840.n64 a_17685_3840.t4 81.437
R1612 a_17685_3840.n31 a_17685_3840.t13 69.653
R1613 a_17685_3840.n32 a_17685_3840.t9 68.683
R1614 a_17685_3840.n63 a_17685_3840.n0 66.545
R1615 a_17685_3840.n62 a_17685_3840.n61 47.861
R1616 a_17685_3840.n24 a_17685_3840.n23 45.936
R1617 a_17685_3840.n32 a_17685_3840.n31 45.7
R1618 a_17685_3840.n30 a_17685_3840.n24 41.108
R1619 a_17685_3840.n61 a_17685_3840.n57 41.07
R1620 a_17685_3840.n65 a_17685_3840.n33 40.118
R1621 a_17685_3840.n0 a_17685_3840.t15 29.277
R1622 a_17685_3840.n0 a_17685_3840.t14 28.576
R1623 a_17685_3840.n0 a_17685_3840.t16 28.565
R1624 a_17685_3840.n33 a_17685_3840.t10 28.565
R1625 a_17685_3840.n33 a_17685_3840.t7 28.565
R1626 a_17685_3840.n67 a_17685_3840.t8 28.565
R1627 a_17685_3840.t11 a_17685_3840.n67 28.565
R1628 a_17685_3840.n56 a_17685_3840.n44 24.999
R1629 a_17685_3840.n65 a_17685_3840.n64 24.605
R1630 a_17685_3840.n23 a_17685_3840.n11 24.399
R1631 a_17685_3840.n34 a_17685_3840.t50 23.529
R1632 a_17685_3840.n1 a_17685_3840.t43 23.485
R1633 a_17685_3840.n12 a_17685_3840.t35 23.474
R1634 a_17685_3840.n45 a_17685_3840.t59 23.456
R1635 a_17685_3840.n66 a_17685_3840.n65 20.217
R1636 a_17685_3840.n66 a_17685_3840.n32 19.791
R1637 a_17685_3840.n44 a_17685_3840.t39 15.401
R1638 a_17685_3840.n11 a_17685_3840.t54 15.374
R1639 a_17685_3840.n55 a_17685_3840.t26 15.341
R1640 a_17685_3840.n22 a_17685_3840.t27 15.334
R1641 a_17685_3840.n23 a_17685_3840.n22 12.228
R1642 a_17685_3840.n56 a_17685_3840.n55 11.433
R1643 a_17685_3840.n43 a_17685_3840.n42 10.674
R1644 a_17685_3840.n42 a_17685_3840.n41 10.674
R1645 a_17685_3840.n41 a_17685_3840.n40 10.674
R1646 a_17685_3840.n40 a_17685_3840.n39 10.674
R1647 a_17685_3840.n39 a_17685_3840.n38 10.674
R1648 a_17685_3840.n38 a_17685_3840.n37 10.674
R1649 a_17685_3840.n37 a_17685_3840.n36 10.674
R1650 a_17685_3840.n36 a_17685_3840.n35 10.674
R1651 a_17685_3840.n35 a_17685_3840.n34 10.674
R1652 a_17685_3840.n21 a_17685_3840.n20 10.655
R1653 a_17685_3840.n20 a_17685_3840.n19 10.655
R1654 a_17685_3840.n19 a_17685_3840.n18 10.655
R1655 a_17685_3840.n18 a_17685_3840.n17 10.655
R1656 a_17685_3840.n17 a_17685_3840.n16 10.655
R1657 a_17685_3840.n16 a_17685_3840.n15 10.655
R1658 a_17685_3840.n15 a_17685_3840.n14 10.655
R1659 a_17685_3840.n14 a_17685_3840.n13 10.655
R1660 a_17685_3840.n13 a_17685_3840.n12 10.655
R1661 a_17685_3840.n10 a_17685_3840.n9 10.637
R1662 a_17685_3840.n9 a_17685_3840.n8 10.637
R1663 a_17685_3840.n8 a_17685_3840.n7 10.637
R1664 a_17685_3840.n7 a_17685_3840.n6 10.637
R1665 a_17685_3840.n6 a_17685_3840.n5 10.637
R1666 a_17685_3840.n5 a_17685_3840.n4 10.637
R1667 a_17685_3840.n4 a_17685_3840.n3 10.637
R1668 a_17685_3840.n3 a_17685_3840.n2 10.637
R1669 a_17685_3840.n2 a_17685_3840.n1 10.637
R1670 a_17685_3840.n54 a_17685_3840.n53 10.625
R1671 a_17685_3840.n53 a_17685_3840.n52 10.625
R1672 a_17685_3840.n52 a_17685_3840.n51 10.625
R1673 a_17685_3840.n51 a_17685_3840.n50 10.625
R1674 a_17685_3840.n50 a_17685_3840.n49 10.625
R1675 a_17685_3840.n49 a_17685_3840.n48 10.625
R1676 a_17685_3840.n48 a_17685_3840.n47 10.625
R1677 a_17685_3840.n47 a_17685_3840.n46 10.625
R1678 a_17685_3840.n46 a_17685_3840.n45 10.625
R1679 a_17685_3840.n45 a_17685_3840.t19 8.716
R1680 a_17685_3840.n46 a_17685_3840.t25 8.716
R1681 a_17685_3840.n47 a_17685_3840.t34 8.716
R1682 a_17685_3840.n48 a_17685_3840.t40 8.716
R1683 a_17685_3840.n49 a_17685_3840.t17 8.716
R1684 a_17685_3840.n50 a_17685_3840.t23 8.716
R1685 a_17685_3840.n51 a_17685_3840.t32 8.716
R1686 a_17685_3840.n52 a_17685_3840.t30 8.716
R1687 a_17685_3840.n53 a_17685_3840.t37 8.716
R1688 a_17685_3840.n54 a_17685_3840.t45 8.716
R1689 a_17685_3840.n1 a_17685_3840.t51 8.713
R1690 a_17685_3840.n2 a_17685_3840.t56 8.713
R1691 a_17685_3840.n3 a_17685_3840.t64 8.713
R1692 a_17685_3840.n4 a_17685_3840.t20 8.713
R1693 a_17685_3840.n5 a_17685_3840.t48 8.713
R1694 a_17685_3840.n6 a_17685_3840.t53 8.713
R1695 a_17685_3840.n7 a_17685_3840.t60 8.713
R1696 a_17685_3840.n8 a_17685_3840.t58 8.713
R1697 a_17685_3840.n9 a_17685_3840.t63 8.713
R1698 a_17685_3840.n10 a_17685_3840.t22 8.713
R1699 a_17685_3840.n12 a_17685_3840.t42 8.708
R1700 a_17685_3840.n13 a_17685_3840.t49 8.708
R1701 a_17685_3840.n14 a_17685_3840.t55 8.708
R1702 a_17685_3840.n15 a_17685_3840.t61 8.708
R1703 a_17685_3840.n16 a_17685_3840.t18 8.708
R1704 a_17685_3840.n17 a_17685_3840.t24 8.708
R1705 a_17685_3840.n18 a_17685_3840.t33 8.708
R1706 a_17685_3840.n19 a_17685_3840.t31 8.708
R1707 a_17685_3840.n20 a_17685_3840.t38 8.708
R1708 a_17685_3840.n21 a_17685_3840.t46 8.708
R1709 a_17685_3840.n43 a_17685_3840.t52 8.704
R1710 a_17685_3840.n34 a_17685_3840.t57 8.704
R1711 a_17685_3840.n35 a_17685_3840.t62 8.704
R1712 a_17685_3840.n36 a_17685_3840.t21 8.704
R1713 a_17685_3840.n37 a_17685_3840.t28 8.704
R1714 a_17685_3840.n38 a_17685_3840.t29 8.704
R1715 a_17685_3840.n39 a_17685_3840.t36 8.704
R1716 a_17685_3840.n40 a_17685_3840.t44 8.704
R1717 a_17685_3840.n41 a_17685_3840.t41 8.704
R1718 a_17685_3840.n42 a_17685_3840.t47 8.704
R1719 a_17685_3840.n22 a_17685_3840.n21 8.14
R1720 a_17685_3840.n44 a_17685_3840.n43 8.128
R1721 a_17685_3840.n55 a_17685_3840.n54 8.116
R1722 a_17685_3840.n11 a_17685_3840.n10 8.112
R1723 a_14266_8900.t16 a_14266_8900.t25 1273.78
R1724 a_14266_8900.n0 a_14266_8900.t47 193.916
R1725 a_14266_8900.t47 a_14266_8900.t53 127.855
R1726 a_14266_8900.t47 a_14266_8900.t21 113.753
R1727 a_14266_8900.t47 a_14266_8900.t11 113.753
R1728 a_14266_8900.t47 a_14266_8900.t32 113.753
R1729 a_14266_8900.t47 a_14266_8900.t41 113.753
R1730 a_14266_8900.t47 a_14266_8900.t52 113.753
R1731 a_14266_8900.t47 a_14266_8900.t50 113.753
R1732 a_14266_8900.t47 a_14266_8900.t58 113.753
R1733 a_14266_8900.t47 a_14266_8900.t18 113.753
R1734 a_14266_8900.t47 a_14266_8900.t8 113.753
R1735 a_14266_8900.t47 a_14266_8900.t48 113.753
R1736 a_14266_8900.t47 a_14266_8900.t42 113.753
R1737 a_14266_8900.t47 a_14266_8900.t54 113.753
R1738 a_14266_8900.t47 a_14266_8900.t17 113.753
R1739 a_14266_8900.t47 a_14266_8900.t34 113.753
R1740 a_14266_8900.t47 a_14266_8900.t45 113.753
R1741 a_14266_8900.t47 a_14266_8900.t39 113.753
R1742 a_14266_8900.t47 a_14266_8900.t13 113.753
R1743 a_14266_8900.t47 a_14266_8900.t5 113.753
R1744 a_14266_8900.t47 a_14266_8900.t29 113.753
R1745 a_14266_8900.t47 a_14266_8900.t23 113.753
R1746 a_14266_8900.t47 a_14266_8900.t51 113.753
R1747 a_14266_8900.t47 a_14266_8900.t59 113.753
R1748 a_14266_8900.t47 a_14266_8900.t20 113.753
R1749 a_14266_8900.t47 a_14266_8900.t9 113.753
R1750 a_14266_8900.t47 a_14266_8900.t49 113.753
R1751 a_14266_8900.t47 a_14266_8900.t43 113.753
R1752 a_14266_8900.t47 a_14266_8900.t55 113.753
R1753 a_14266_8900.t47 a_14266_8900.t19 113.753
R1754 a_14266_8900.t47 a_14266_8900.t35 113.753
R1755 a_14266_8900.t47 a_14266_8900.t46 113.753
R1756 a_14266_8900.t47 a_14266_8900.t40 113.753
R1757 a_14266_8900.t47 a_14266_8900.t14 113.753
R1758 a_14266_8900.t47 a_14266_8900.t6 113.753
R1759 a_14266_8900.t47 a_14266_8900.t30 113.753
R1760 a_14266_8900.t47 a_14266_8900.t24 113.753
R1761 a_14266_8900.t47 a_14266_8900.t2 113.753
R1762 a_14266_8900.t47 a_14266_8900.t60 113.753
R1763 a_14266_8900.t47 a_14266_8900.t27 113.753
R1764 a_14266_8900.t47 a_14266_8900.t36 113.753
R1765 a_14266_8900.t47 a_14266_8900.t31 113.753
R1766 a_14266_8900.t47 a_14266_8900.t57 113.753
R1767 a_14266_8900.t47 a_14266_8900.t56 113.753
R1768 a_14266_8900.t47 a_14266_8900.t7 113.753
R1769 a_14266_8900.t47 a_14266_8900.t22 113.753
R1770 a_14266_8900.t47 a_14266_8900.t15 113.753
R1771 a_14266_8900.t47 a_14266_8900.t33 113.753
R1772 a_14266_8900.t47 a_14266_8900.t44 113.753
R1773 a_14266_8900.t47 a_14266_8900.t38 113.753
R1774 a_14266_8900.t47 a_14266_8900.t12 113.753
R1775 a_14266_8900.t47 a_14266_8900.t4 113.753
R1776 a_14266_8900.t47 a_14266_8900.t28 113.753
R1777 a_14266_8900.t47 a_14266_8900.t37 113.753
R1778 a_14266_8900.t47 a_14266_8900.t10 113.753
R1779 a_14266_8900.t47 a_14266_8900.t3 113.753
R1780 a_14266_8900.t47 a_14266_8900.t26 113.753
R1781 a_14266_8900.t1 a_14266_8900.t16 57.619
R1782 a_14266_8900.t16 a_14266_8900.n0 53.144
R1783 a_14266_8900.n0 a_14266_8900.t0 28.571
R1784 a_22629_11500.n6 a_22629_11500.n4 75.711
R1785 a_22629_11500.n1 a_22629_11500.n0 75.707
R1786 a_22629_11500.n2 a_22629_11500.n1 75.707
R1787 a_22629_11500.n3 a_22629_11500.n2 75.707
R1788 a_22629_11500.n4 a_22629_11500.n3 75.707
R1789 a_22629_11500.n0 a_22629_11500.n5 75.707
R1790 a_22629_11500.n4 a_22629_11500.t11 17.401
R1791 a_22629_11500.n3 a_22629_11500.t13 17.401
R1792 a_22629_11500.n2 a_22629_11500.t8 17.401
R1793 a_22629_11500.n1 a_22629_11500.t10 17.401
R1794 a_22629_11500.n0 a_22629_11500.t9 17.401
R1795 a_22629_11500.n4 a_22629_11500.t2 17.4
R1796 a_22629_11500.n3 a_22629_11500.t0 17.4
R1797 a_22629_11500.n2 a_22629_11500.t3 17.4
R1798 a_22629_11500.n1 a_22629_11500.t1 17.4
R1799 a_22629_11500.n0 a_22629_11500.t4 17.4
R1800 a_22629_11500.n5 a_22629_11500.t7 17.4
R1801 a_22629_11500.n5 a_22629_11500.t5 17.4
R1802 a_22629_11500.n6 a_22629_11500.t12 17.4
R1803 a_22629_11500.t6 a_22629_11500.n6 17.4
R1804 a_66357_25280.t0 a_66357_25280.t1 87.142
R1805 a_63529_26290.n1 a_63529_26290.t5 350.253
R1806 a_63529_26290.n1 a_63529_26290.t4 189.586
R1807 a_63529_26290.n2 a_63529_26290.n1 97.205
R1808 a_63529_26290.n3 a_63529_26290.t0 89.119
R1809 a_63529_26290.n2 a_63529_26290.n0 79.305
R1810 a_63529_26290.n3 a_63529_26290.n2 66.705
R1811 a_63529_26290.n0 a_63529_26290.t2 63.333
R1812 a_63529_26290.t1 a_63529_26290.n3 41.041
R1813 a_63529_26290.n0 a_63529_26290.t3 31.979
R1814 a_63419_26414.t0 a_63419_26414.n0 194.654
R1815 a_63419_26414.n0 a_63419_26414.t1 168.384
R1816 a_63419_26414.n0 a_63419_26414.t2 63.321
R1817 a_28478_5597.n0 a_28478_5597.n1 75.71
R1818 a_28478_5597.n4 a_28478_5597.n5 75.708
R1819 a_28478_5597.n2 a_28478_5597.n3 75.707
R1820 a_28478_5597.n3 a_28478_5597.n4 75.707
R1821 a_28478_5597.n1 a_28478_5597.n6 75.707
R1822 a_28478_5597.n0 a_28478_5597.n2 75.706
R1823 a_28478_5597.t8 a_28478_5597.n0 17.401
R1824 a_28478_5597.n4 a_28478_5597.t2 17.401
R1825 a_28478_5597.n3 a_28478_5597.t7 17.401
R1826 a_28478_5597.n2 a_28478_5597.t3 17.401
R1827 a_28478_5597.n1 a_28478_5597.t6 17.401
R1828 a_28478_5597.n5 a_28478_5597.t5 17.4
R1829 a_28478_5597.n5 a_28478_5597.t12 17.4
R1830 a_28478_5597.n4 a_28478_5597.t11 17.4
R1831 a_28478_5597.n3 a_28478_5597.t0 17.4
R1832 a_28478_5597.n2 a_28478_5597.t9 17.4
R1833 a_28478_5597.n1 a_28478_5597.t13 17.4
R1834 a_28478_5597.n6 a_28478_5597.t4 17.4
R1835 a_28478_5597.n6 a_28478_5597.t10 17.4
R1836 a_28478_5597.n0 a_28478_5597.t1 17.4
R1837 a_29252_5597.n0 a_29252_5597.n6 75.709
R1838 a_29252_5597.n4 a_29252_5597.n5 75.708
R1839 a_29252_5597.n1 a_29252_5597.n2 75.707
R1840 a_29252_5597.n2 a_29252_5597.n3 75.707
R1841 a_29252_5597.n3 a_29252_5597.n4 75.707
R1842 a_29252_5597.n0 a_29252_5597.n1 75.706
R1843 a_29252_5597.n0 a_29252_5597.t13 17.401
R1844 a_29252_5597.n4 a_29252_5597.t0 17.401
R1845 a_29252_5597.n3 a_29252_5597.t4 17.401
R1846 a_29252_5597.n2 a_29252_5597.t1 17.401
R1847 a_29252_5597.n1 a_29252_5597.t5 17.401
R1848 a_29252_5597.n5 a_29252_5597.t3 17.4
R1849 a_29252_5597.n5 a_29252_5597.t11 17.4
R1850 a_29252_5597.n4 a_29252_5597.t8 17.4
R1851 a_29252_5597.n3 a_29252_5597.t6 17.4
R1852 a_29252_5597.n2 a_29252_5597.t9 17.4
R1853 a_29252_5597.n1 a_29252_5597.t7 17.4
R1854 a_29252_5597.n6 a_29252_5597.t2 17.4
R1855 a_29252_5597.n6 a_29252_5597.t10 17.4
R1856 a_29252_5597.t12 a_29252_5597.n0 17.4
R1857 a_29510_5597.n6 a_29510_5597.n4 75.711
R1858 a_29510_5597.n1 a_29510_5597.n0 75.707
R1859 a_29510_5597.n2 a_29510_5597.n1 75.707
R1860 a_29510_5597.n3 a_29510_5597.n2 75.707
R1861 a_29510_5597.n4 a_29510_5597.n3 75.707
R1862 a_29510_5597.n0 a_29510_5597.n5 75.707
R1863 a_29510_5597.n4 a_29510_5597.t4 17.401
R1864 a_29510_5597.n3 a_29510_5597.t0 17.401
R1865 a_29510_5597.n2 a_29510_5597.t5 17.401
R1866 a_29510_5597.n1 a_29510_5597.t1 17.401
R1867 a_29510_5597.n0 a_29510_5597.t6 17.401
R1868 a_29510_5597.n4 a_29510_5597.t9 17.4
R1869 a_29510_5597.n3 a_29510_5597.t7 17.4
R1870 a_29510_5597.n2 a_29510_5597.t10 17.4
R1871 a_29510_5597.n1 a_29510_5597.t8 17.4
R1872 a_29510_5597.n0 a_29510_5597.t13 17.4
R1873 a_29510_5597.n5 a_29510_5597.t2 17.4
R1874 a_29510_5597.n5 a_29510_5597.t11 17.4
R1875 a_29510_5597.n6 a_29510_5597.t3 17.4
R1876 a_29510_5597.t12 a_29510_5597.n6 17.4
R1877 Vso3b.n0 Vso3b.t1 17.996
R1878 Vso3b Vso3b.n0 0.383
R1879 Vso3b Vso3b.n1 6.01
R1880 Vso3b.n1 Vso3b.t4 412.212
R1881 Vso3b.n1 Vso3b.n3 141.4
R1882 Vso3b.n3 Vso3b.t5 289.757
R1883 Vso3b.n3 Vso3b.n2 63.152
R1884 Vso3b.n2 Vso3b.t2 375.287
R1885 Vso3b.n2 Vso3b.t3 391.653
R1886 Vso3b.n0 Vso3b.t0 132.37
R1887 a_8744_13422.t0 a_8744_13422.t1 53.512
R1888 Vso5b.n0 Vso5b.t1 17.996
R1889 Vso5b.n1 Vso5b.n0 0.455
R1890 Vso5b Vso5b.n1 0.127
R1891 Vso5b.n1 Vso5b.n2 2.498
R1892 Vso5b.n2 Vso5b.t4 413.786
R1893 Vso5b.n2 Vso5b.n4 138.132
R1894 Vso5b.n4 Vso5b.t5 291.452
R1895 Vso5b.n4 Vso5b.n3 59.644
R1896 Vso5b.n3 Vso5b.t2 378.337
R1897 Vso5b.n3 Vso5b.t3 388.603
R1898 Vso5b.n0 Vso5b.t0 132.37
R1899 a_8748_12270.t0 a_8748_12270.t1 53.512
R1900 a_23661_5596.n0 a_23661_5596.n3 75.71
R1901 a_23661_5596.n4 a_23661_5596.n5 75.708
R1902 a_23661_5596.n2 a_23661_5596.n1 75.707
R1903 a_23661_5596.n3 a_23661_5596.n2 75.707
R1904 a_23661_5596.n1 a_23661_5596.n6 75.707
R1905 a_23661_5596.n0 a_23661_5596.n4 75.706
R1906 a_23661_5596.n0 a_23661_5596.t8 17.401
R1907 a_23661_5596.n4 a_23661_5596.t10 17.401
R1908 a_23661_5596.n3 a_23661_5596.t11 17.401
R1909 a_23661_5596.n2 a_23661_5596.t9 17.401
R1910 a_23661_5596.n1 a_23661_5596.t7 17.401
R1911 a_23661_5596.n5 a_23661_5596.t13 17.4
R1912 a_23661_5596.n5 a_23661_5596.t4 17.4
R1913 a_23661_5596.n4 a_23661_5596.t1 17.4
R1914 a_23661_5596.n3 a_23661_5596.t2 17.4
R1915 a_23661_5596.n2 a_23661_5596.t0 17.4
R1916 a_23661_5596.n1 a_23661_5596.t5 17.4
R1917 a_23661_5596.n6 a_23661_5596.t12 17.4
R1918 a_23661_5596.n6 a_23661_5596.t3 17.4
R1919 a_23661_5596.t6 a_23661_5596.n0 17.4
R1920 a_52052_20860.t0 a_52052_20860.n16 2527.24
R1921 a_52052_20860.n8 a_52052_20860.t6 212.622
R1922 a_52052_20860.n5 a_52052_20860.t18 212.622
R1923 a_52052_20860.n12 a_52052_20860.n10 208.271
R1924 a_52052_20860.n2 a_52052_20860.n0 208.271
R1925 a_52052_20860.n14 a_52052_20860.n12 208.271
R1926 a_52052_20860.n9 a_52052_20860.n8 208.271
R1927 a_52052_20860.n4 a_52052_20860.n2 208.271
R1928 a_52052_20860.n6 a_52052_20860.n5 208.271
R1929 a_52052_20860.n7 a_52052_20860.n6 122.265
R1930 a_52052_20860.n15 a_52052_20860.n14 121.297
R1931 a_52052_20860.n7 a_52052_20860.n4 63.478
R1932 a_52052_20860.n15 a_52052_20860.n9 63.217
R1933 a_52052_20860.n16 a_52052_20860.n7 38.746
R1934 a_52052_20860.n16 a_52052_20860.n15 15.694
R1935 a_52052_20860.n8 a_52052_20860.t8 4.351
R1936 a_52052_20860.n9 a_52052_20860.t4 4.351
R1937 a_52052_20860.n5 a_52052_20860.t15 4.351
R1938 a_52052_20860.n6 a_52052_20860.t12 4.351
R1939 a_52052_20860.n10 a_52052_20860.t9 4.35
R1940 a_52052_20860.n10 a_52052_20860.t5 4.35
R1941 a_52052_20860.n11 a_52052_20860.t7 4.35
R1942 a_52052_20860.n11 a_52052_20860.t1 4.35
R1943 a_52052_20860.n13 a_52052_20860.t2 4.35
R1944 a_52052_20860.n13 a_52052_20860.t3 4.35
R1945 a_52052_20860.n0 a_52052_20860.t16 4.35
R1946 a_52052_20860.n0 a_52052_20860.t17 4.35
R1947 a_52052_20860.n1 a_52052_20860.t10 4.35
R1948 a_52052_20860.n1 a_52052_20860.t13 4.35
R1949 a_52052_20860.n3 a_52052_20860.t14 4.35
R1950 a_52052_20860.n3 a_52052_20860.t11 4.35
R1951 a_52052_20860.n14 a_52052_20860.n13 0.001
R1952 a_52052_20860.n12 a_52052_20860.n11 0.001
R1953 a_52052_20860.n4 a_52052_20860.n3 0.001
R1954 a_52052_20860.n2 a_52052_20860.n1 0.001
R1955 a_56334_20860.t0 a_56334_20860.n0 171.567
R1956 a_56334_20860.n0 a_56334_20860.t1 171.564
R1957 a_56334_20860.n0 a_56334_20860.t2 171.52
R1958 a_23156_5032.n0 a_23156_5032.t7 365.308
R1959 a_23156_5032.n4 a_23156_5032.t2 93.107
R1960 a_23156_5032.n5 a_23156_5032.n4 75.71
R1961 a_23156_5032.n3 a_23156_5032.n2 75.707
R1962 a_23156_5032.n2 a_23156_5032.n1 75.707
R1963 a_23156_5032.n1 a_23156_5032.n0 75.707
R1964 a_23156_5032.n5 a_23156_5032.n3 75.706
R1965 a_23156_5032.t6 a_23156_5032.n5 17.401
R1966 a_23156_5032.n0 a_23156_5032.t3 17.401
R1967 a_23156_5032.n1 a_23156_5032.t0 17.401
R1968 a_23156_5032.n2 a_23156_5032.t5 17.401
R1969 a_23156_5032.n3 a_23156_5032.t1 17.401
R1970 a_23156_5032.n4 a_23156_5032.t4 17.401
R1971 a_28478_17218.n0 a_28478_17218.n2 75.71
R1972 a_28478_17218.n4 a_28478_17218.n5 75.708
R1973 a_28478_17218.n2 a_28478_17218.n1 75.707
R1974 a_28478_17218.n3 a_28478_17218.n4 75.707
R1975 a_28478_17218.n1 a_28478_17218.n6 75.707
R1976 a_28478_17218.n0 a_28478_17218.n3 75.706
R1977 a_28478_17218.t6 a_28478_17218.n0 17.401
R1978 a_28478_17218.n4 a_28478_17218.t5 17.401
R1979 a_28478_17218.n3 a_28478_17218.t2 17.401
R1980 a_28478_17218.n2 a_28478_17218.t3 17.401
R1981 a_28478_17218.n1 a_28478_17218.t4 17.401
R1982 a_28478_17218.n5 a_28478_17218.t1 17.4
R1983 a_28478_17218.n5 a_28478_17218.t10 17.4
R1984 a_28478_17218.n4 a_28478_17218.t7 17.4
R1985 a_28478_17218.n3 a_28478_17218.t11 17.4
R1986 a_28478_17218.n2 a_28478_17218.t12 17.4
R1987 a_28478_17218.n1 a_28478_17218.t13 17.4
R1988 a_28478_17218.n6 a_28478_17218.t0 17.4
R1989 a_28478_17218.n6 a_28478_17218.t9 17.4
R1990 a_28478_17218.n0 a_28478_17218.t8 17.4
R1991 a_65546_25646.n0 a_65546_25646.t1 194.654
R1992 a_65546_25646.t0 a_65546_25646.n0 168.384
R1993 a_65546_25646.n0 a_65546_25646.t2 63.321
R1994 a_23436_16644.t12 a_23436_16644.t43 1273.78
R1995 a_23436_16644.n0 a_23436_16644.t1 1158.7
R1996 a_23436_16644.n0 a_23436_16644.t12 169.095
R1997 a_23436_16644.t12 a_23436_16644.t53 134.91
R1998 a_23436_16644.t12 a_23436_16644.t45 113.753
R1999 a_23436_16644.t12 a_23436_16644.t5 113.753
R2000 a_23436_16644.t12 a_23436_16644.t21 113.753
R2001 a_23436_16644.t12 a_23436_16644.t20 113.753
R2002 a_23436_16644.t12 a_23436_16644.t2 113.753
R2003 a_23436_16644.t12 a_23436_16644.t17 113.753
R2004 a_23436_16644.t12 a_23436_16644.t37 113.753
R2005 a_23436_16644.t12 a_23436_16644.t33 113.753
R2006 a_23436_16644.t12 a_23436_16644.t44 113.753
R2007 a_23436_16644.t12 a_23436_16644.t58 113.753
R2008 a_23436_16644.t12 a_23436_16644.t14 113.753
R2009 a_23436_16644.t12 a_23436_16644.t32 113.753
R2010 a_23436_16644.t12 a_23436_16644.t10 113.753
R2011 a_23436_16644.t12 a_23436_16644.t28 113.753
R2012 a_23436_16644.t12 a_23436_16644.t26 113.753
R2013 a_23436_16644.t12 a_23436_16644.t34 113.753
R2014 a_23436_16644.t12 a_23436_16644.t46 113.753
R2015 a_23436_16644.t12 a_23436_16644.t6 113.753
R2016 a_23436_16644.t12 a_23436_16644.t24 113.753
R2017 a_23436_16644.t12 a_23436_16644.t49 113.753
R2018 a_23436_16644.t12 a_23436_16644.t22 113.753
R2019 a_23436_16644.t12 a_23436_16644.t40 113.753
R2020 a_23436_16644.t12 a_23436_16644.t57 113.753
R2021 a_23436_16644.t12 a_23436_16644.t55 113.753
R2022 a_23436_16644.t12 a_23436_16644.t8 113.753
R2023 a_23436_16644.t12 a_23436_16644.t18 113.753
R2024 a_23436_16644.t12 a_23436_16644.t38 113.753
R2025 a_23436_16644.t12 a_23436_16644.t11 113.753
R2026 a_23436_16644.t12 a_23436_16644.t29 113.753
R2027 a_23436_16644.t12 a_23436_16644.t27 113.753
R2028 a_23436_16644.t12 a_23436_16644.t35 113.753
R2029 a_23436_16644.t12 a_23436_16644.t47 113.753
R2030 a_23436_16644.t12 a_23436_16644.t7 113.753
R2031 a_23436_16644.t12 a_23436_16644.t25 113.753
R2032 a_23436_16644.t12 a_23436_16644.t50 113.753
R2033 a_23436_16644.t12 a_23436_16644.t23 113.753
R2034 a_23436_16644.t12 a_23436_16644.t41 113.753
R2035 a_23436_16644.t12 a_23436_16644.t59 113.753
R2036 a_23436_16644.t12 a_23436_16644.t56 113.753
R2037 a_23436_16644.t12 a_23436_16644.t9 113.753
R2038 a_23436_16644.t12 a_23436_16644.t19 113.753
R2039 a_23436_16644.t12 a_23436_16644.t39 113.753
R2040 a_23436_16644.t12 a_23436_16644.t54 113.753
R2041 a_23436_16644.t12 a_23436_16644.t15 113.753
R2042 a_23436_16644.t12 a_23436_16644.t36 113.753
R2043 a_23436_16644.t12 a_23436_16644.t52 113.753
R2044 a_23436_16644.t12 a_23436_16644.t51 113.753
R2045 a_23436_16644.t12 a_23436_16644.t4 113.753
R2046 a_23436_16644.t12 a_23436_16644.t13 113.753
R2047 a_23436_16644.t12 a_23436_16644.t31 113.753
R2048 a_23436_16644.t12 a_23436_16644.t48 113.753
R2049 a_23436_16644.t12 a_23436_16644.t30 113.753
R2050 a_23436_16644.t12 a_23436_16644.t42 113.753
R2051 a_23436_16644.t12 a_23436_16644.t3 113.753
R2052 a_23436_16644.t12 a_23436_16644.t16 113.753
R2053 a_23436_16644.t0 a_23436_16644.n0 59.624
R2054 a_25299_17217.n0 a_25299_17217.n1 75.71
R2055 a_25299_17217.n4 a_25299_17217.n5 75.708
R2056 a_25299_17217.n2 a_25299_17217.n3 75.707
R2057 a_25299_17217.n3 a_25299_17217.n4 75.707
R2058 a_25299_17217.n1 a_25299_17217.n6 75.707
R2059 a_25299_17217.n0 a_25299_17217.n2 75.706
R2060 a_25299_17217.n0 a_25299_17217.t11 17.401
R2061 a_25299_17217.n4 a_25299_17217.t8 17.401
R2062 a_25299_17217.n3 a_25299_17217.t13 17.401
R2063 a_25299_17217.n2 a_25299_17217.t9 17.401
R2064 a_25299_17217.n1 a_25299_17217.t10 17.401
R2065 a_25299_17217.n5 a_25299_17217.t12 17.4
R2066 a_25299_17217.n5 a_25299_17217.t3 17.4
R2067 a_25299_17217.n4 a_25299_17217.t0 17.4
R2068 a_25299_17217.n3 a_25299_17217.t4 17.4
R2069 a_25299_17217.n2 a_25299_17217.t1 17.4
R2070 a_25299_17217.n1 a_25299_17217.t5 17.4
R2071 a_25299_17217.n6 a_25299_17217.t7 17.4
R2072 a_25299_17217.n6 a_25299_17217.t2 17.4
R2073 a_25299_17217.t6 a_25299_17217.n0 17.4
R2074 a_26589_17217.n0 a_26589_17217.n4 75.71
R2075 a_26589_17217.n2 a_26589_17217.n1 75.707
R2076 a_26589_17217.n3 a_26589_17217.n2 75.707
R2077 a_26589_17217.n4 a_26589_17217.n3 75.707
R2078 a_26589_17217.n1 a_26589_17217.n6 75.707
R2079 a_26589_17217.n0 a_26589_17217.n5 75.707
R2080 a_26589_17217.t0 a_26589_17217.n0 17.401
R2081 a_26589_17217.n4 a_26589_17217.t3 17.401
R2082 a_26589_17217.n3 a_26589_17217.t1 17.401
R2083 a_26589_17217.n2 a_26589_17217.t9 17.401
R2084 a_26589_17217.n1 a_26589_17217.t8 17.401
R2085 a_26589_17217.n5 a_26589_17217.t2 17.4
R2086 a_26589_17217.n5 a_26589_17217.t10 17.4
R2087 a_26589_17217.n4 a_26589_17217.t11 17.4
R2088 a_26589_17217.n3 a_26589_17217.t4 17.4
R2089 a_26589_17217.n2 a_26589_17217.t12 17.4
R2090 a_26589_17217.n1 a_26589_17217.t6 17.4
R2091 a_26589_17217.n6 a_26589_17217.t7 17.4
R2092 a_26589_17217.n6 a_26589_17217.t5 17.4
R2093 a_26589_17217.n0 a_26589_17217.t13 17.4
R2094 a_26847_17217.n4 a_26847_17217.n5 75.708
R2095 a_26847_17217.n0 a_26847_17217.n1 75.707
R2096 a_26847_17217.n1 a_26847_17217.n2 75.707
R2097 a_26847_17217.n2 a_26847_17217.n3 75.707
R2098 a_26847_17217.n3 a_26847_17217.n4 75.707
R2099 a_26847_17217.n6 a_26847_17217.n0 75.707
R2100 a_26847_17217.n4 a_26847_17217.t13 17.401
R2101 a_26847_17217.n3 a_26847_17217.t0 17.401
R2102 a_26847_17217.n2 a_26847_17217.t11 17.401
R2103 a_26847_17217.n1 a_26847_17217.t12 17.401
R2104 a_26847_17217.n0 a_26847_17217.t1 17.401
R2105 a_26847_17217.n5 a_26847_17217.t10 17.4
R2106 a_26847_17217.n5 a_26847_17217.t3 17.4
R2107 a_26847_17217.n4 a_26847_17217.t7 17.4
R2108 a_26847_17217.n3 a_26847_17217.t4 17.4
R2109 a_26847_17217.n2 a_26847_17217.t8 17.4
R2110 a_26847_17217.n1 a_26847_17217.t6 17.4
R2111 a_26847_17217.n0 a_26847_17217.t5 17.4
R2112 a_26847_17217.n6 a_26847_17217.t2 17.4
R2113 a_26847_17217.t9 a_26847_17217.n6 17.4
R2114 a_51636_13108.t0 a_51636_13108.n0 14.331
R2115 a_51636_13108.n0 a_51636_13108.n3 3.54
R2116 a_51636_13108.n3 a_51636_13108.n11 8.062
R2117 a_51636_13108.n10 a_51636_13108.t6 96.508
R2118 a_51636_13108.n11 a_51636_13108.n10 0.138
R2119 a_51636_13108.n5 a_51636_13108.t9 96.486
R2120 a_51636_13108.n9 a_51636_13108.t12 96.489
R2121 a_51636_13108.n5 a_51636_13108.n9 0.667
R2122 a_51636_13108.n7 a_51636_13108.n5 0.002
R2123 a_51636_13108.n10 a_51636_13108.n7 0.646
R2124 a_51636_13108.n8 a_51636_13108.t8 96.96
R2125 a_51636_13108.n8 a_51636_13108.t11 96.486
R2126 a_51636_13108.n9 a_51636_13108.n8 0.286
R2127 a_51636_13108.n6 a_51636_13108.t13 96.96
R2128 a_51636_13108.n6 a_51636_13108.t7 96.486
R2129 a_51636_13108.n7 a_51636_13108.n6 0.286
R2130 a_51636_13108.n4 a_51636_13108.t10 96.96
R2131 a_51636_13108.n4 a_51636_13108.t5 96.486
R2132 a_51636_13108.n11 a_51636_13108.n4 0.3
R2133 a_51636_13108.n3 a_51636_13108.t4 607.174
R2134 a_51636_13108.n1 a_51636_13108.n2 4.438
R2135 a_51636_13108.n0 a_51636_13108.n1 3.405
R2136 a_51636_13108.n2 a_51636_13108.t1 17.451
R2137 a_51636_13108.n2 a_51636_13108.t2 17.452
R2138 a_51636_13108.n1 a_51636_13108.t3 14.302
R2139 a_51276_14152.t1 a_51276_14152.n0 14.331
R2140 a_51276_14152.n0 a_51276_14152.n1 0.394
R2141 a_51276_14152.n7 a_51276_14152.t0 17.453
R2142 a_51276_14152.n0 a_51276_14152.n7 2.815
R2143 a_51276_14152.n7 a_51276_14152.t3 17.451
R2144 a_51276_14152.n1 a_51276_14152.t2 14.505
R2145 a_51276_14152.n1 a_51276_14152.n6 227.496
R2146 a_51276_14152.n3 a_51276_14152.n4 0.003
R2147 a_51276_14152.n6 a_51276_14152.n3 48.522
R2148 a_51276_14152.n3 a_51276_14152.n5 153.01
R2149 a_51276_14152.n5 a_51276_14152.t5 8.7
R2150 a_51276_14152.n5 a_51276_14152.t8 8.7
R2151 a_51276_14152.n4 a_51276_14152.t9 8.7
R2152 a_51276_14152.n4 a_51276_14152.t4 8.7
R2153 a_51276_14152.n6 a_51276_14152.n2 123.385
R2154 a_51276_14152.n2 a_51276_14152.t7 153.199
R2155 a_51276_14152.n2 a_51276_14152.t6 8.703
R2156 a_25557_5596.n6 a_25557_5596.n4 75.44
R2157 a_25557_5596.n1 a_25557_5596.n0 75.436
R2158 a_25557_5596.n2 a_25557_5596.n1 75.436
R2159 a_25557_5596.n3 a_25557_5596.n2 75.436
R2160 a_25557_5596.n4 a_25557_5596.n3 75.436
R2161 a_25557_5596.n0 a_25557_5596.n5 75.436
R2162 a_25557_5596.n4 a_25557_5596.t5 17.401
R2163 a_25557_5596.n3 a_25557_5596.t6 17.401
R2164 a_25557_5596.n2 a_25557_5596.t2 17.401
R2165 a_25557_5596.n1 a_25557_5596.t4 17.401
R2166 a_25557_5596.n0 a_25557_5596.t1 17.401
R2167 a_25557_5596.n4 a_25557_5596.t8 17.4
R2168 a_25557_5596.n3 a_25557_5596.t13 17.4
R2169 a_25557_5596.n2 a_25557_5596.t11 17.4
R2170 a_25557_5596.n1 a_25557_5596.t7 17.4
R2171 a_25557_5596.n0 a_25557_5596.t10 17.4
R2172 a_25557_5596.n5 a_25557_5596.t3 17.4
R2173 a_25557_5596.n5 a_25557_5596.t12 17.4
R2174 a_25557_5596.t0 a_25557_5596.n6 17.4
R2175 a_25557_5596.n6 a_25557_5596.t9 17.4
R2176 a_25815_5596.n0 a_25815_5596.n6 75.709
R2177 a_25815_5596.n4 a_25815_5596.n5 75.708
R2178 a_25815_5596.n1 a_25815_5596.n2 75.707
R2179 a_25815_5596.n2 a_25815_5596.n3 75.707
R2180 a_25815_5596.n3 a_25815_5596.n4 75.707
R2181 a_25815_5596.n0 a_25815_5596.n1 75.706
R2182 a_25815_5596.n0 a_25815_5596.t0 17.401
R2183 a_25815_5596.n4 a_25815_5596.t9 17.401
R2184 a_25815_5596.n3 a_25815_5596.t1 17.401
R2185 a_25815_5596.n2 a_25815_5596.t10 17.401
R2186 a_25815_5596.n1 a_25815_5596.t11 17.401
R2187 a_25815_5596.n5 a_25815_5596.t13 17.4
R2188 a_25815_5596.n5 a_25815_5596.t7 17.4
R2189 a_25815_5596.n4 a_25815_5596.t4 17.4
R2190 a_25815_5596.n3 a_25815_5596.t2 17.4
R2191 a_25815_5596.n2 a_25815_5596.t5 17.4
R2192 a_25815_5596.n1 a_25815_5596.t3 17.4
R2193 a_25815_5596.n6 a_25815_5596.t12 17.4
R2194 a_25815_5596.n6 a_25815_5596.t6 17.4
R2195 a_25815_5596.t8 a_25815_5596.n0 17.4
R2196 a_62795_26048.n3 a_62795_26048.t5 530.008
R2197 a_62795_26048.n2 a_62795_26048.t6 334.888
R2198 a_62795_26048.n7 a_62795_26048.t3 255.459
R2199 a_62795_26048.n5 a_62795_26048.t4 224.611
R2200 a_62795_26048.n2 a_62795_26048.t7 196.882
R2201 a_62795_26048.n3 a_62795_26048.t2 141.921
R2202 a_62795_26048.t0 a_62795_26048.n8 126.03
R2203 a_62795_26048.n0 a_62795_26048.t1 99.672
R2204 a_62795_26048.n4 a_62795_26048.n3 92.562
R2205 a_62795_26048.n4 a_62795_26048.n2 44.57
R2206 a_62795_26048.n0 a_62795_26048.n4 38.638
R2207 a_62795_26048.n1 a_62795_26048.n6 15
R2208 a_62795_26048.n8 a_62795_26048.n7 15
R2209 a_62795_26048.n1 a_62795_26048.n5 13.653
R2210 a_62795_26048.n8 a_62795_26048.n1 3.182
R2211 a_62795_26048.n1 a_62795_26048.n0 2.692
R2212 a_63216_26048.n1 a_63216_26048.n0 163.71
R2213 a_63216_26048.t1 a_63216_26048.n1 82.083
R2214 a_63216_26048.n0 a_63216_26048.t0 63.333
R2215 a_63216_26048.n1 a_63216_26048.t2 63.321
R2216 a_63216_26048.n0 a_63216_26048.t3 29.726
R2217 a_63311_26048.n1 a_63311_26048.t5 332.579
R2218 a_63311_26048.n1 a_63311_26048.t4 168.699
R2219 a_63311_26048.n2 a_63311_26048.n1 104.381
R2220 a_63311_26048.n2 a_63311_26048.n0 101.869
R2221 a_63311_26048.t1 a_63311_26048.n3 96.154
R2222 a_63311_26048.n3 a_63311_26048.n2 92.648
R2223 a_63311_26048.n3 a_63311_26048.t2 65.666
R2224 a_63311_26048.n0 a_63311_26048.t0 65
R2225 a_63311_26048.n0 a_63311_26048.t3 45
R2226 a_26073_11500.n0 a_26073_11500.n6 75.709
R2227 a_26073_11500.n4 a_26073_11500.n5 75.708
R2228 a_26073_11500.n1 a_26073_11500.n2 75.707
R2229 a_26073_11500.n2 a_26073_11500.n3 75.707
R2230 a_26073_11500.n3 a_26073_11500.n4 75.707
R2231 a_26073_11500.n0 a_26073_11500.n1 75.706
R2232 a_26073_11500.t0 a_26073_11500.n0 17.401
R2233 a_26073_11500.n4 a_26073_11500.t6 17.401
R2234 a_26073_11500.n3 a_26073_11500.t1 17.401
R2235 a_26073_11500.n2 a_26073_11500.t13 17.401
R2236 a_26073_11500.n1 a_26073_11500.t2 17.401
R2237 a_26073_11500.n5 a_26073_11500.t4 17.4
R2238 a_26073_11500.n5 a_26073_11500.t5 17.4
R2239 a_26073_11500.n4 a_26073_11500.t8 17.4
R2240 a_26073_11500.n3 a_26073_11500.t11 17.4
R2241 a_26073_11500.n2 a_26073_11500.t9 17.4
R2242 a_26073_11500.n1 a_26073_11500.t10 17.4
R2243 a_26073_11500.n6 a_26073_11500.t3 17.4
R2244 a_26073_11500.n6 a_26073_11500.t12 17.4
R2245 a_26073_11500.n0 a_26073_11500.t7 17.4
R2246 a_26331_11500.n0 a_26331_11500.n1 75.71
R2247 a_26331_11500.n4 a_26331_11500.n5 75.708
R2248 a_26331_11500.n2 a_26331_11500.n3 75.707
R2249 a_26331_11500.n3 a_26331_11500.n4 75.707
R2250 a_26331_11500.n1 a_26331_11500.n6 75.707
R2251 a_26331_11500.n0 a_26331_11500.n2 75.706
R2252 a_26331_11500.n0 a_26331_11500.t13 17.401
R2253 a_26331_11500.n4 a_26331_11500.t7 17.401
R2254 a_26331_11500.n3 a_26331_11500.t12 17.401
R2255 a_26331_11500.n2 a_26331_11500.t8 17.401
R2256 a_26331_11500.n1 a_26331_11500.t9 17.401
R2257 a_26331_11500.n5 a_26331_11500.t11 17.4
R2258 a_26331_11500.n5 a_26331_11500.t4 17.4
R2259 a_26331_11500.n4 a_26331_11500.t0 17.4
R2260 a_26331_11500.n3 a_26331_11500.t5 17.4
R2261 a_26331_11500.n2 a_26331_11500.t1 17.4
R2262 a_26331_11500.n1 a_26331_11500.t2 17.4
R2263 a_26331_11500.n6 a_26331_11500.t10 17.4
R2264 a_26331_11500.n6 a_26331_11500.t3 17.4
R2265 a_26331_11500.t6 a_26331_11500.n0 17.4
R2266 a_28220_5597.n0 a_28220_5597.n1 75.439
R2267 a_28220_5597.n4 a_28220_5597.n5 75.437
R2268 a_28220_5597.n2 a_28220_5597.n3 75.436
R2269 a_28220_5597.n3 a_28220_5597.n4 75.436
R2270 a_28220_5597.n1 a_28220_5597.n6 75.436
R2271 a_28220_5597.n0 a_28220_5597.n2 75.435
R2272 a_28220_5597.t11 a_28220_5597.n0 17.401
R2273 a_28220_5597.n4 a_28220_5597.t5 17.401
R2274 a_28220_5597.n3 a_28220_5597.t10 17.401
R2275 a_28220_5597.n2 a_28220_5597.t6 17.401
R2276 a_28220_5597.n1 a_28220_5597.t9 17.401
R2277 a_28220_5597.n5 a_28220_5597.t8 17.4
R2278 a_28220_5597.n5 a_28220_5597.t3 17.4
R2279 a_28220_5597.n4 a_28220_5597.t0 17.4
R2280 a_28220_5597.n3 a_28220_5597.t12 17.4
R2281 a_28220_5597.n2 a_28220_5597.t1 17.4
R2282 a_28220_5597.n1 a_28220_5597.t4 17.4
R2283 a_28220_5597.n6 a_28220_5597.t7 17.4
R2284 a_28220_5597.n6 a_28220_5597.t2 17.4
R2285 a_28220_5597.n0 a_28220_5597.t13 17.4
R2286 CLK_IN.n0 CLK_IN.t1 17.996
R2287 CLK_IN.n1 CLK_IN.n0 1.608
R2288 CLK_IN CLK_IN.n5 10.221
R2289 CLK_IN CLK_IN.n1 64.808
R2290 CLK_IN.n5 CLK_IN.t5 211.008
R2291 CLK_IN.n5 CLK_IN.t4 294.554
R2292 CLK_IN.n1 CLK_IN.n4 7.694
R2293 CLK_IN.n4 CLK_IN.t3 423.069
R2294 CLK_IN.n4 CLK_IN.n3 155.549
R2295 CLK_IN.n3 CLK_IN.t6 292.807
R2296 CLK_IN.n3 CLK_IN.n2 56.933
R2297 CLK_IN.n2 CLK_IN.t7 378.337
R2298 CLK_IN.n2 CLK_IN.t2 388.603
R2299 CLK_IN.n0 CLK_IN.t0 132.37
R2300 a_4288_11534.t1 a_4288_11534.n0 17.028
R2301 a_4288_11534.n0 a_4288_11534.t2 18.871
R2302 a_4288_11534.n0 a_4288_11534.n1 1.817
R2303 a_4288_11534.n1 a_4288_11534.n2 5.932
R2304 a_4288_11534.n2 a_4288_11534.t3 597.139
R2305 a_4288_11534.n2 a_4288_11534.t4 434.044
R2306 a_4288_11534.n1 a_4288_11534.t0 26.804
R2307 a_26847_5596.n0 a_26847_5596.n1 75.71
R2308 a_26847_5596.n4 a_26847_5596.n5 75.708
R2309 a_26847_5596.n2 a_26847_5596.n3 75.707
R2310 a_26847_5596.n3 a_26847_5596.n4 75.707
R2311 a_26847_5596.n1 a_26847_5596.n6 75.707
R2312 a_26847_5596.n0 a_26847_5596.n2 75.706
R2313 a_26847_5596.n0 a_26847_5596.t2 17.401
R2314 a_26847_5596.n4 a_26847_5596.t9 17.401
R2315 a_26847_5596.n3 a_26847_5596.t1 17.401
R2316 a_26847_5596.n2 a_26847_5596.t3 17.401
R2317 a_26847_5596.n1 a_26847_5596.t8 17.401
R2318 a_26847_5596.n5 a_26847_5596.t7 17.4
R2319 a_26847_5596.n5 a_26847_5596.t11 17.4
R2320 a_26847_5596.n4 a_26847_5596.t5 17.4
R2321 a_26847_5596.n3 a_26847_5596.t13 17.4
R2322 a_26847_5596.n2 a_26847_5596.t6 17.4
R2323 a_26847_5596.n1 a_26847_5596.t12 17.4
R2324 a_26847_5596.n6 a_26847_5596.t4 17.4
R2325 a_26847_5596.n6 a_26847_5596.t10 17.4
R2326 a_26847_5596.t0 a_26847_5596.n0 17.4
R2327 a_25778_4988.n0 a_25778_4988.t0 334.707
R2328 a_25778_4988.n2 a_25778_4988.t3 93.107
R2329 a_25778_4988.n5 a_25778_4988.n4 75.71
R2330 a_25778_4988.n3 a_25778_4988.n2 75.707
R2331 a_25778_4988.n4 a_25778_4988.n3 75.707
R2332 a_25778_4988.n1 a_25778_4988.n0 75.707
R2333 a_25778_4988.n5 a_25778_4988.n1 75.706
R2334 a_25778_4988.t6 a_25778_4988.n5 17.401
R2335 a_25778_4988.n0 a_25778_4988.t4 17.401
R2336 a_25778_4988.n1 a_25778_4988.t1 17.401
R2337 a_25778_4988.n4 a_25778_4988.t2 17.401
R2338 a_25778_4988.n3 a_25778_4988.t7 17.401
R2339 a_25778_4988.n2 a_25778_4988.t5 17.401
R2340 Fvco.t0 Fvco.n0 77.367
R2341 Fvco.n0 Fvco.t1 28.578
R2342 Fvco.n81 Fvco.n0 132.569
R2343 Fvco.n80 Fvco.n81 0.428
R2344 Fvco Fvco.n80 0.038
R2345 Fvco.n80 Fvco.n79 1.398
R2346 Fvco.n79 Fvco.t11 1273.78
R2347 Fvco.n79 Fvco.t34 1.21
R2348 Fvco.n81 Fvco.n1 3.526
R2349 Fvco.n2 Fvco.t23 113.753
R2350 Fvco.n3 Fvco.t4 113.753
R2351 Fvco.n4 Fvco.t6 113.753
R2352 Fvco.n5 Fvco.t37 113.753
R2353 Fvco.n1 Fvco.n5 0.175
R2354 Fvco.n5 Fvco.n4 0.325
R2355 Fvco.n4 Fvco.n3 0.325
R2356 Fvco.n3 Fvco.n2 0.325
R2357 Fvco.n2 Fvco.n6 0.522
R2358 Fvco.n7 Fvco.t56 113.753
R2359 Fvco.n8 Fvco.t38 113.753
R2360 Fvco.n9 Fvco.t42 113.753
R2361 Fvco.n10 Fvco.t5 113.753
R2362 Fvco.n11 Fvco.t8 113.753
R2363 Fvco.n12 Fvco.t61 113.753
R2364 Fvco.n13 Fvco.t43 113.753
R2365 Fvco.n14 Fvco.t49 113.753
R2366 Fvco.n78 Fvco.n14 0.158
R2367 Fvco.n14 Fvco.n13 0.168
R2368 Fvco.n13 Fvco.n12 0.168
R2369 Fvco.n12 Fvco.n11 0.168
R2370 Fvco.n9 Fvco.n10 0.168
R2371 Fvco.n8 Fvco.n9 0.168
R2372 Fvco.n7 Fvco.n8 0.168
R2373 Fvco.n6 Fvco.n7 0.21
R2374 Fvco.n22 Fvco.n23 0.32
R2375 Fvco.n21 Fvco.n22 0.328
R2376 Fvco.n20 Fvco.n21 0.32
R2377 Fvco.n19 Fvco.n20 0.335
R2378 Fvco.n78 Fvco.n19 0.32
R2379 Fvco.n23 Fvco.n26 0.536
R2380 Fvco.n26 Fvco.n25 0.248
R2381 Fvco.n28 Fvco.n24 0.211
R2382 Fvco.n77 Fvco.n28 0.005
R2383 Fvco.n27 Fvco.n77 0.085
R2384 Fvco.n77 Fvco.t32 0.145
R2385 Fvco.n31 Fvco.n27 0.206
R2386 Fvco.n30 Fvco.n31 0.248
R2387 Fvco.n29 Fvco.n30 0.248
R2388 Fvco.n32 Fvco.n29 0.462
R2389 Fvco.n33 Fvco.t60 113.753
R2390 Fvco.n34 Fvco.t46 113.753
R2391 Fvco.n35 Fvco.t51 113.753
R2392 Fvco.n36 Fvco.t14 113.753
R2393 Fvco.n37 Fvco.t20 113.753
R2394 Fvco.n38 Fvco.t3 113.753
R2395 Fvco.n39 Fvco.t53 113.753
R2396 Fvco.n40 Fvco.t55 113.753
R2397 Fvco.n23 Fvco.n40 0.158
R2398 Fvco.n40 Fvco.n39 0.168
R2399 Fvco.n37 Fvco.n38 0.168
R2400 Fvco.n36 Fvco.n37 0.168
R2401 Fvco.n35 Fvco.n36 0.168
R2402 Fvco.n34 Fvco.n35 0.168
R2403 Fvco.n33 Fvco.n34 0.168
R2404 Fvco.n32 Fvco.n33 0.21
R2405 Fvco.n41 Fvco.t22 113.753
R2406 Fvco.n42 Fvco.t26 113.753
R2407 Fvco.n43 Fvco.t10 113.753
R2408 Fvco.n44 Fvco.t16 113.753
R2409 Fvco.n45 Fvco.t41 113.753
R2410 Fvco.n46 Fvco.t48 113.753
R2411 Fvco.n47 Fvco.t35 113.753
R2412 Fvco.n48 Fvco.t18 113.753
R2413 Fvco.n22 Fvco.n41 0.158
R2414 Fvco.n41 Fvco.n48 0.168
R2415 Fvco.n46 Fvco.n47 0.168
R2416 Fvco.n45 Fvco.n46 0.168
R2417 Fvco.n44 Fvco.n45 0.168
R2418 Fvco.n43 Fvco.n44 0.168
R2419 Fvco.n42 Fvco.n43 0.168
R2420 Fvco.n76 Fvco.n42 0.21
R2421 Fvco.n76 Fvco.n32 0.171
R2422 Fvco.n49 Fvco.n76 0.178
R2423 Fvco.n50 Fvco.t59 113.753
R2424 Fvco.n51 Fvco.t45 113.753
R2425 Fvco.n52 Fvco.t50 113.753
R2426 Fvco.n53 Fvco.t12 113.753
R2427 Fvco.n54 Fvco.t19 113.753
R2428 Fvco.n55 Fvco.t2 113.753
R2429 Fvco.n56 Fvco.t52 113.753
R2430 Fvco.n57 Fvco.t54 113.753
R2431 Fvco.n21 Fvco.n57 0.158
R2432 Fvco.n57 Fvco.n56 0.168
R2433 Fvco.n56 Fvco.n55 0.168
R2434 Fvco.n53 Fvco.n54 0.168
R2435 Fvco.n52 Fvco.n53 0.168
R2436 Fvco.n51 Fvco.n52 0.168
R2437 Fvco.n50 Fvco.n51 0.168
R2438 Fvco.n49 Fvco.n50 0.21
R2439 Fvco.n58 Fvco.t21 113.753
R2440 Fvco.n59 Fvco.t25 113.753
R2441 Fvco.n60 Fvco.t9 113.753
R2442 Fvco.n61 Fvco.t15 113.753
R2443 Fvco.n62 Fvco.t40 113.753
R2444 Fvco.n63 Fvco.t47 113.753
R2445 Fvco.n64 Fvco.t33 113.753
R2446 Fvco.n65 Fvco.t17 113.753
R2447 Fvco.n20 Fvco.n58 0.158
R2448 Fvco.n58 Fvco.n65 0.168
R2449 Fvco.n65 Fvco.n64 0.168
R2450 Fvco.n62 Fvco.n63 0.168
R2451 Fvco.n61 Fvco.n62 0.168
R2452 Fvco.n60 Fvco.n61 0.168
R2453 Fvco.n59 Fvco.n60 0.168
R2454 Fvco.n75 Fvco.n59 0.21
R2455 Fvco.n75 Fvco.n49 0.171
R2456 Fvco.n66 Fvco.n75 0.186
R2457 Fvco.n67 Fvco.t36 113.753
R2458 Fvco.n68 Fvco.t24 113.753
R2459 Fvco.n69 Fvco.t27 113.753
R2460 Fvco.n70 Fvco.t57 113.753
R2461 Fvco.n71 Fvco.t58 113.753
R2462 Fvco.n72 Fvco.t44 113.753
R2463 Fvco.n73 Fvco.t28 113.753
R2464 Fvco.n74 Fvco.t30 113.753
R2465 Fvco.n19 Fvco.n74 0.158
R2466 Fvco.n74 Fvco.n73 0.168
R2467 Fvco.n73 Fvco.n72 0.168
R2468 Fvco.n72 Fvco.n71 0.168
R2469 Fvco.n69 Fvco.n70 0.168
R2470 Fvco.n68 Fvco.n69 0.168
R2471 Fvco.n67 Fvco.n68 0.168
R2472 Fvco.n66 Fvco.n67 0.21
R2473 Fvco.n6 Fvco.n66 0.171
R2474 Fvco.n15 Fvco.t39 113.753
R2475 Fvco.n16 Fvco.t31 113.753
R2476 Fvco.n17 Fvco.t7 113.753
R2477 Fvco.n18 Fvco.t13 113.753
R2478 Fvco.n18 Fvco.n78 0.597
R2479 Fvco.n17 Fvco.n18 0.325
R2480 Fvco.n16 Fvco.n17 0.325
R2481 Fvco.n15 Fvco.n16 0.325
R2482 Fvco.n1 Fvco.n15 0.102
R2483 Fvco.n1 Fvco.t29 0.4
R2484 a_22887_17217.n0 a_22887_17217.n6 75.438
R2485 a_22887_17217.n4 a_22887_17217.n5 75.437
R2486 a_22887_17217.n1 a_22887_17217.n2 75.436
R2487 a_22887_17217.n2 a_22887_17217.n3 75.436
R2488 a_22887_17217.n3 a_22887_17217.n4 75.436
R2489 a_22887_17217.n0 a_22887_17217.n1 75.435
R2490 a_22887_17217.n0 a_22887_17217.t6 17.401
R2491 a_22887_17217.n4 a_22887_17217.t3 17.401
R2492 a_22887_17217.n3 a_22887_17217.t13 17.401
R2493 a_22887_17217.n2 a_22887_17217.t4 17.401
R2494 a_22887_17217.n1 a_22887_17217.t7 17.401
R2495 a_22887_17217.n5 a_22887_17217.t11 17.4
R2496 a_22887_17217.n5 a_22887_17217.t12 17.4
R2497 a_22887_17217.n4 a_22887_17217.t9 17.4
R2498 a_22887_17217.n3 a_22887_17217.t5 17.4
R2499 a_22887_17217.n2 a_22887_17217.t8 17.4
R2500 a_22887_17217.n1 a_22887_17217.t1 17.4
R2501 a_22887_17217.n6 a_22887_17217.t10 17.4
R2502 a_22887_17217.n6 a_22887_17217.t2 17.4
R2503 a_22887_17217.t0 a_22887_17217.n0 17.4
R2504 a_23145_17217.n0 a_23145_17217.n3 75.71
R2505 a_23145_17217.n4 a_23145_17217.n5 75.708
R2506 a_23145_17217.n2 a_23145_17217.n1 75.707
R2507 a_23145_17217.n3 a_23145_17217.n2 75.707
R2508 a_23145_17217.n1 a_23145_17217.n6 75.707
R2509 a_23145_17217.n0 a_23145_17217.n4 75.706
R2510 a_23145_17217.n0 a_23145_17217.t7 17.401
R2511 a_23145_17217.n4 a_23145_17217.t11 17.401
R2512 a_23145_17217.n3 a_23145_17217.t12 17.401
R2513 a_23145_17217.n2 a_23145_17217.t13 17.401
R2514 a_23145_17217.n1 a_23145_17217.t8 17.401
R2515 a_23145_17217.n5 a_23145_17217.t10 17.4
R2516 a_23145_17217.n5 a_23145_17217.t5 17.4
R2517 a_23145_17217.n4 a_23145_17217.t2 17.4
R2518 a_23145_17217.n3 a_23145_17217.t3 17.4
R2519 a_23145_17217.n2 a_23145_17217.t1 17.4
R2520 a_23145_17217.n1 a_23145_17217.t0 17.4
R2521 a_23145_17217.n6 a_23145_17217.t9 17.4
R2522 a_23145_17217.n6 a_23145_17217.t4 17.4
R2523 a_23145_17217.t6 a_23145_17217.n0 17.4
R2524 a_56602_11692.t1 a_56602_11692.n0 14.474
R2525 a_56602_11692.n0 a_56602_11692.n10 0.497
R2526 a_56602_11692.n11 a_56602_11692.t0 17.453
R2527 a_56602_11692.n10 a_56602_11692.n11 1.13
R2528 a_56602_11692.n11 a_56602_11692.t3 17.451
R2529 a_56602_11692.n10 a_56602_11692.n1 886.086
R2530 a_56602_11692.n1 a_56602_11692.n9 446.23
R2531 a_56602_11692.n7 a_56602_11692.t9 212.622
R2532 a_56602_11692.n8 a_56602_11692.n7 208.271
R2533 a_56602_11692.n9 a_56602_11692.n8 73.665
R2534 a_56602_11692.n8 a_56602_11692.t7 4.351
R2535 a_56602_11692.n7 a_56602_11692.t4 4.351
R2536 a_56602_11692.n3 a_56602_11692.n4 0.001
R2537 a_56602_11692.n5 a_56602_11692.n6 0.001
R2538 a_56602_11692.n3 a_56602_11692.n2 208.271
R2539 a_56602_11692.n5 a_56602_11692.n3 208.271
R2540 a_56602_11692.n9 a_56602_11692.n5 164.114
R2541 a_56602_11692.n6 a_56602_11692.t11 4.35
R2542 a_56602_11692.n6 a_56602_11692.t12 4.35
R2543 a_56602_11692.n4 a_56602_11692.t8 4.35
R2544 a_56602_11692.n4 a_56602_11692.t10 4.35
R2545 a_56602_11692.n2 a_56602_11692.t5 4.35
R2546 a_56602_11692.n2 a_56602_11692.t6 4.35
R2547 a_56602_11692.n1 a_56602_11692.t13 5.714
R2548 a_56602_11692.n0 a_56602_11692.t2 14.302
R2549 vbiasob.n0 vbiasob.t0 67.964
R2550 vbiasob vbiasob.t3 61.399
R2551 vbiasob vbiasob.t4 60.299
R2552 vbiasob.n0 vbiasob.t2 18.573
R2553 vbiasob vbiasob.n0 13.139
R2554 vbiasob.n0 vbiasob.t1 6.729
R2555 a_56272_15934.t1 a_56272_15934.t0 409.924
R2556 a_27962_5597.n0 a_27962_5597.n3 75.71
R2557 a_27962_5597.n4 a_27962_5597.n5 75.708
R2558 a_27962_5597.n2 a_27962_5597.n1 75.707
R2559 a_27962_5597.n3 a_27962_5597.n2 75.707
R2560 a_27962_5597.n1 a_27962_5597.n6 75.707
R2561 a_27962_5597.n0 a_27962_5597.n4 75.706
R2562 a_27962_5597.n0 a_27962_5597.t12 17.401
R2563 a_27962_5597.n4 a_27962_5597.t7 17.401
R2564 a_27962_5597.n3 a_27962_5597.t8 17.401
R2565 a_27962_5597.n2 a_27962_5597.t13 17.401
R2566 a_27962_5597.n1 a_27962_5597.t11 17.401
R2567 a_27962_5597.n5 a_27962_5597.t10 17.4
R2568 a_27962_5597.n5 a_27962_5597.t4 17.4
R2569 a_27962_5597.n4 a_27962_5597.t1 17.4
R2570 a_27962_5597.n3 a_27962_5597.t2 17.4
R2571 a_27962_5597.n2 a_27962_5597.t0 17.4
R2572 a_27962_5597.n1 a_27962_5597.t5 17.4
R2573 a_27962_5597.n6 a_27962_5597.t9 17.4
R2574 a_27962_5597.n6 a_27962_5597.t3 17.4
R2575 a_27962_5597.t6 a_27962_5597.n0 17.4
R2576 a_54966_2992.t0 a_54966_2992.t1 25.776
R2577 vbiasbuffer.n0 vbiasbuffer.t0 136.915
R2578 vbiasbuffer vbiasbuffer.t4 125.304
R2579 vbiasbuffer vbiasbuffer.t3 120.586
R2580 vbiasbuffer.n0 vbiasbuffer.t2 22.405
R2581 vbiasbuffer vbiasbuffer.n0 15.641
R2582 vbiasbuffer.n0 vbiasbuffer.t1 5.719
R2583 a_26073_17217.n0 a_26073_17217.n1 75.71
R2584 a_26073_17217.n4 a_26073_17217.n5 75.708
R2585 a_26073_17217.n2 a_26073_17217.n3 75.707
R2586 a_26073_17217.n3 a_26073_17217.n4 75.707
R2587 a_26073_17217.n1 a_26073_17217.n6 75.707
R2588 a_26073_17217.n0 a_26073_17217.n2 75.706
R2589 a_26073_17217.n0 a_26073_17217.t13 17.401
R2590 a_26073_17217.n4 a_26073_17217.t9 17.401
R2591 a_26073_17217.n3 a_26073_17217.t6 17.401
R2592 a_26073_17217.n2 a_26073_17217.t10 17.401
R2593 a_26073_17217.n1 a_26073_17217.t7 17.401
R2594 a_26073_17217.n5 a_26073_17217.t12 17.4
R2595 a_26073_17217.n5 a_26073_17217.t3 17.4
R2596 a_26073_17217.n4 a_26073_17217.t8 17.4
R2597 a_26073_17217.n3 a_26073_17217.t5 17.4
R2598 a_26073_17217.n2 a_26073_17217.t4 17.4
R2599 a_26073_17217.n1 a_26073_17217.t2 17.4
R2600 a_26073_17217.n6 a_26073_17217.t11 17.4
R2601 a_26073_17217.n6 a_26073_17217.t1 17.4
R2602 a_26073_17217.t0 a_26073_17217.n0 17.4
R2603 a_26331_17217.n0 a_26331_17217.n6 75.709
R2604 a_26331_17217.n4 a_26331_17217.n5 75.708
R2605 a_26331_17217.n1 a_26331_17217.n2 75.707
R2606 a_26331_17217.n2 a_26331_17217.n3 75.707
R2607 a_26331_17217.n3 a_26331_17217.n4 75.707
R2608 a_26331_17217.n0 a_26331_17217.n1 75.706
R2609 a_26331_17217.n0 a_26331_17217.t13 17.401
R2610 a_26331_17217.n4 a_26331_17217.t8 17.401
R2611 a_26331_17217.n3 a_26331_17217.t12 17.401
R2612 a_26331_17217.n2 a_26331_17217.t9 17.401
R2613 a_26331_17217.n1 a_26331_17217.t7 17.401
R2614 a_26331_17217.n5 a_26331_17217.t11 17.4
R2615 a_26331_17217.n5 a_26331_17217.t4 17.4
R2616 a_26331_17217.n4 a_26331_17217.t1 17.4
R2617 a_26331_17217.n3 a_26331_17217.t5 17.4
R2618 a_26331_17217.n2 a_26331_17217.t2 17.4
R2619 a_26331_17217.n1 a_26331_17217.t0 17.4
R2620 a_26331_17217.n6 a_26331_17217.t10 17.4
R2621 a_26331_17217.n6 a_26331_17217.t3 17.4
R2622 a_26331_17217.t6 a_26331_17217.n0 17.4
R2623 a_57726_5786.n0 a_57726_5786.t3 85.561
R2624 a_57726_5786.n0 a_57726_5786.t1 85.561
R2625 a_57726_5786.n0 a_57726_5786.t5 39.685
R2626 a_57726_5786.n0 a_57726_5786.t0 17.517
R2627 a_57726_5786.t4 a_57726_5786.n0 6.973
R2628 a_57726_5786.n0 a_57726_5786.t2 5.8
R2629 a_25299_11500.n0 a_25299_11500.n1 75.71
R2630 a_25299_11500.n4 a_25299_11500.n5 75.708
R2631 a_25299_11500.n2 a_25299_11500.n3 75.707
R2632 a_25299_11500.n3 a_25299_11500.n4 75.707
R2633 a_25299_11500.n1 a_25299_11500.n6 75.707
R2634 a_25299_11500.n0 a_25299_11500.n2 75.706
R2635 a_25299_11500.n0 a_25299_11500.t8 17.401
R2636 a_25299_11500.n4 a_25299_11500.t10 17.401
R2637 a_25299_11500.n3 a_25299_11500.t7 17.401
R2638 a_25299_11500.n2 a_25299_11500.t11 17.401
R2639 a_25299_11500.n1 a_25299_11500.t12 17.401
R2640 a_25299_11500.n5 a_25299_11500.t9 17.4
R2641 a_25299_11500.n5 a_25299_11500.t4 17.4
R2642 a_25299_11500.n4 a_25299_11500.t0 17.4
R2643 a_25299_11500.n3 a_25299_11500.t5 17.4
R2644 a_25299_11500.n2 a_25299_11500.t1 17.4
R2645 a_25299_11500.n1 a_25299_11500.t2 17.4
R2646 a_25299_11500.n6 a_25299_11500.t13 17.4
R2647 a_25299_11500.n6 a_25299_11500.t3 17.4
R2648 a_25299_11500.t6 a_25299_11500.n0 17.4
R2649 a_25557_11500.n4 a_25557_11500.n5 75.437
R2650 a_25557_11500.n0 a_25557_11500.n1 75.436
R2651 a_25557_11500.n1 a_25557_11500.n2 75.436
R2652 a_25557_11500.n2 a_25557_11500.n3 75.436
R2653 a_25557_11500.n3 a_25557_11500.n4 75.436
R2654 a_25557_11500.n6 a_25557_11500.n0 75.436
R2655 a_25557_11500.n4 a_25557_11500.t1 17.401
R2656 a_25557_11500.n3 a_25557_11500.t3 17.401
R2657 a_25557_11500.n2 a_25557_11500.t5 17.401
R2658 a_25557_11500.n1 a_25557_11500.t0 17.401
R2659 a_25557_11500.n0 a_25557_11500.t2 17.401
R2660 a_25557_11500.n5 a_25557_11500.t4 17.4
R2661 a_25557_11500.n5 a_25557_11500.t6 17.4
R2662 a_25557_11500.n4 a_25557_11500.t9 17.4
R2663 a_25557_11500.n3 a_25557_11500.t7 17.4
R2664 a_25557_11500.n2 a_25557_11500.t10 17.4
R2665 a_25557_11500.n1 a_25557_11500.t8 17.4
R2666 a_25557_11500.n0 a_25557_11500.t11 17.4
R2667 a_25557_11500.n6 a_25557_11500.t13 17.4
R2668 a_25557_11500.t12 a_25557_11500.n6 17.4
R2669 a_25299_5596.n0 a_25299_5596.n6 75.709
R2670 a_25299_5596.n4 a_25299_5596.n5 75.708
R2671 a_25299_5596.n1 a_25299_5596.n2 75.707
R2672 a_25299_5596.n2 a_25299_5596.n3 75.707
R2673 a_25299_5596.n3 a_25299_5596.n4 75.707
R2674 a_25299_5596.n0 a_25299_5596.n1 75.706
R2675 a_25299_5596.n0 a_25299_5596.t13 17.401
R2676 a_25299_5596.n4 a_25299_5596.t9 17.401
R2677 a_25299_5596.n3 a_25299_5596.t7 17.401
R2678 a_25299_5596.n2 a_25299_5596.t10 17.401
R2679 a_25299_5596.n1 a_25299_5596.t8 17.401
R2680 a_25299_5596.n5 a_25299_5596.t12 17.4
R2681 a_25299_5596.n5 a_25299_5596.t5 17.4
R2682 a_25299_5596.n4 a_25299_5596.t2 17.4
R2683 a_25299_5596.n3 a_25299_5596.t0 17.4
R2684 a_25299_5596.n2 a_25299_5596.t3 17.4
R2685 a_25299_5596.n1 a_25299_5596.t1 17.4
R2686 a_25299_5596.n6 a_25299_5596.t11 17.4
R2687 a_25299_5596.n6 a_25299_5596.t4 17.4
R2688 a_25299_5596.t6 a_25299_5596.n0 17.4
R2689 a_26589_5596.n0 a_26589_5596.n3 75.71
R2690 a_26589_5596.n4 a_26589_5596.n5 75.708
R2691 a_26589_5596.n2 a_26589_5596.n1 75.707
R2692 a_26589_5596.n3 a_26589_5596.n2 75.707
R2693 a_26589_5596.n1 a_26589_5596.n6 75.707
R2694 a_26589_5596.n0 a_26589_5596.n4 75.706
R2695 a_26589_5596.t12 a_26589_5596.n0 17.401
R2696 a_26589_5596.n4 a_26589_5596.t7 17.401
R2697 a_26589_5596.n3 a_26589_5596.t8 17.401
R2698 a_26589_5596.n2 a_26589_5596.t13 17.401
R2699 a_26589_5596.n1 a_26589_5596.t11 17.401
R2700 a_26589_5596.n5 a_26589_5596.t10 17.4
R2701 a_26589_5596.n5 a_26589_5596.t4 17.4
R2702 a_26589_5596.n4 a_26589_5596.t5 17.4
R2703 a_26589_5596.n3 a_26589_5596.t6 17.4
R2704 a_26589_5596.n2 a_26589_5596.t0 17.4
R2705 a_26589_5596.n1 a_26589_5596.t1 17.4
R2706 a_26589_5596.n6 a_26589_5596.t9 17.4
R2707 a_26589_5596.n6 a_26589_5596.t3 17.4
R2708 a_26589_5596.n0 a_26589_5596.t2 17.4
R2709 a_28578_5014.n0 a_28578_5014.t0 265.845
R2710 a_28578_5014.t6 a_28578_5014.n5 93.107
R2711 a_28578_5014.n5 a_28578_5014.n4 75.707
R2712 a_28578_5014.n4 a_28578_5014.n3 75.707
R2713 a_28578_5014.n3 a_28578_5014.n2 75.707
R2714 a_28578_5014.n2 a_28578_5014.n1 75.707
R2715 a_28578_5014.n1 a_28578_5014.n0 75.707
R2716 a_28578_5014.n0 a_28578_5014.t7 17.401
R2717 a_28578_5014.n1 a_28578_5014.t4 17.401
R2718 a_28578_5014.n2 a_28578_5014.t2 17.401
R2719 a_28578_5014.n3 a_28578_5014.t5 17.401
R2720 a_28578_5014.n4 a_28578_5014.t3 17.401
R2721 a_28578_5014.n5 a_28578_5014.t1 17.401
R2722 a_23919_11500.n0 a_23919_11500.n4 75.71
R2723 a_23919_11500.n2 a_23919_11500.n1 75.707
R2724 a_23919_11500.n3 a_23919_11500.n2 75.707
R2725 a_23919_11500.n4 a_23919_11500.n3 75.707
R2726 a_23919_11500.n1 a_23919_11500.n6 75.707
R2727 a_23919_11500.n0 a_23919_11500.n5 75.707
R2728 a_23919_11500.t0 a_23919_11500.n0 17.401
R2729 a_23919_11500.n4 a_23919_11500.t2 17.401
R2730 a_23919_11500.n3 a_23919_11500.t1 17.401
R2731 a_23919_11500.n2 a_23919_11500.t3 17.401
R2732 a_23919_11500.n1 a_23919_11500.t5 17.401
R2733 a_23919_11500.n5 a_23919_11500.t4 17.4
R2734 a_23919_11500.n5 a_23919_11500.t9 17.4
R2735 a_23919_11500.n4 a_23919_11500.t10 17.4
R2736 a_23919_11500.n3 a_23919_11500.t12 17.4
R2737 a_23919_11500.n2 a_23919_11500.t7 17.4
R2738 a_23919_11500.n1 a_23919_11500.t13 17.4
R2739 a_23919_11500.n6 a_23919_11500.t6 17.4
R2740 a_23919_11500.n6 a_23919_11500.t11 17.4
R2741 a_23919_11500.n0 a_23919_11500.t8 17.4
R2742 a_24177_11500.n4 a_24177_11500.n5 75.708
R2743 a_24177_11500.n0 a_24177_11500.n1 75.707
R2744 a_24177_11500.n1 a_24177_11500.n2 75.707
R2745 a_24177_11500.n2 a_24177_11500.n3 75.707
R2746 a_24177_11500.n3 a_24177_11500.n4 75.707
R2747 a_24177_11500.n6 a_24177_11500.n0 75.707
R2748 a_24177_11500.n4 a_24177_11500.t10 17.401
R2749 a_24177_11500.n3 a_24177_11500.t12 17.401
R2750 a_24177_11500.n2 a_24177_11500.t11 17.401
R2751 a_24177_11500.n1 a_24177_11500.t13 17.401
R2752 a_24177_11500.n0 a_24177_11500.t8 17.401
R2753 a_24177_11500.n5 a_24177_11500.t7 17.4
R2754 a_24177_11500.n5 a_24177_11500.t0 17.4
R2755 a_24177_11500.n4 a_24177_11500.t3 17.4
R2756 a_24177_11500.n3 a_24177_11500.t1 17.4
R2757 a_24177_11500.n2 a_24177_11500.t4 17.4
R2758 a_24177_11500.n1 a_24177_11500.t2 17.4
R2759 a_24177_11500.n0 a_24177_11500.t5 17.4
R2760 a_24177_11500.n6 a_24177_11500.t9 17.4
R2761 a_24177_11500.t6 a_24177_11500.n6 17.4
R2762 a_50583_13108.n0 a_50583_13108.t0 1776.66
R2763 a_50583_13108.n0 a_50583_13108.t2 171.607
R2764 a_50583_13108.t1 a_50583_13108.n0 171.607
R2765 a_51041_13108.t1 a_51041_13108.n9 15.976
R2766 a_51041_13108.n10 a_51041_13108.n11 1.885
R2767 a_51041_13108.n9 a_51041_13108.n10 3.23
R2768 a_51041_13108.n11 a_51041_13108.t3 18.036
R2769 a_51041_13108.n11 a_51041_13108.t0 17.538
R2770 a_51041_13108.n10 a_51041_13108.t2 14.302
R2771 a_51041_13108.n9 a_51041_13108.n0 741.937
R2772 a_51041_13108.n0 a_51041_13108.n8 362.558
R2773 a_51041_13108.n7 a_51041_13108.t6 96.497
R2774 a_51041_13108.n8 a_51041_13108.n7 0.132
R2775 a_51041_13108.n2 a_51041_13108.t9 96.486
R2776 a_51041_13108.n6 a_51041_13108.t12 96.492
R2777 a_51041_13108.n2 a_51041_13108.n6 0.665
R2778 a_51041_13108.n4 a_51041_13108.n2 0.004
R2779 a_51041_13108.n7 a_51041_13108.n4 0.643
R2780 a_51041_13108.n5 a_51041_13108.t8 96.96
R2781 a_51041_13108.n5 a_51041_13108.t11 96.486
R2782 a_51041_13108.n6 a_51041_13108.n5 0.294
R2783 a_51041_13108.n3 a_51041_13108.t13 96.96
R2784 a_51041_13108.n3 a_51041_13108.t7 96.486
R2785 a_51041_13108.n4 a_51041_13108.n3 0.294
R2786 a_51041_13108.n1 a_51041_13108.t10 96.96
R2787 a_51041_13108.n1 a_51041_13108.t5 96.486
R2788 a_51041_13108.n8 a_51041_13108.n1 0.263
R2789 a_51041_13108.n0 a_51041_13108.t4 930.639
R2790 a_27762_11446.t11 a_27762_11446.t47 1273.78
R2791 a_27762_11446.t11 a_27762_11446.t13 113.753
R2792 a_27762_11446.t11 a_27762_11446.t23 113.753
R2793 a_27762_11446.t11 a_27762_11446.t39 113.753
R2794 a_27762_11446.t11 a_27762_11446.t55 113.753
R2795 a_27762_11446.t11 a_27762_11446.t45 113.753
R2796 a_27762_11446.t11 a_27762_11446.t59 113.753
R2797 a_27762_11446.t11 a_27762_11446.t9 113.753
R2798 a_27762_11446.t11 a_27762_11446.t30 113.753
R2799 a_27762_11446.t21 a_27762_11446.t25 113.753
R2800 a_27762_11446.t21 a_27762_11446.t37 113.753
R2801 a_27762_11446.t21 a_27762_11446.t52 113.753
R2802 a_27762_11446.t21 a_27762_11446.t7 113.753
R2803 a_27762_11446.t11 a_27762_11446.t28 113.753
R2804 a_27762_11446.t11 a_27762_11446.t41 113.753
R2805 a_27762_11446.t21 a_27762_11446.t57 113.753
R2806 a_27762_11446.t21 a_27762_11446.t50 113.753
R2807 a_27762_11446.t21 a_27762_11446.t5 113.753
R2808 a_27762_11446.t21 a_27762_11446.t20 113.753
R2809 a_27762_11446.t21 a_27762_11446.t35 113.753
R2810 a_27762_11446.t11 a_27762_11446.t15 113.753
R2811 a_27762_11446.t11 a_27762_11446.t46 113.753
R2812 a_27762_11446.t11 a_27762_11446.t60 113.753
R2813 a_27762_11446.t11 a_27762_11446.t10 113.753
R2814 a_27762_11446.t21 a_27762_11446.t31 113.753
R2815 a_27762_11446.t21 a_27762_11446.t26 113.753
R2816 a_27762_11446.t21 a_27762_11446.t38 113.753
R2817 a_27762_11446.t21 a_27762_11446.t53 113.753
R2818 a_27762_11446.t21 a_27762_11446.t8 113.753
R2819 a_27762_11446.t11 a_27762_11446.t29 113.753
R2820 a_27762_11446.t21 a_27762_11446.t42 113.753
R2821 a_27762_11446.t21 a_27762_11446.t58 113.753
R2822 a_27762_11446.t21 a_27762_11446.t51 113.753
R2823 a_27762_11446.t21 a_27762_11446.t6 113.753
R2824 a_27762_11446.t21 a_27762_11446.t22 113.753
R2825 a_27762_11446.t21 a_27762_11446.t36 113.753
R2826 a_27762_11446.t11 a_27762_11446.t16 113.753
R2827 a_27762_11446.t11 a_27762_11446.t3 113.753
R2828 a_27762_11446.t11 a_27762_11446.t17 113.753
R2829 a_27762_11446.t21 a_27762_11446.t32 113.753
R2830 a_27762_11446.t21 a_27762_11446.t44 113.753
R2831 a_27762_11446.t21 a_27762_11446.t43 113.753
R2832 a_27762_11446.t21 a_27762_11446.t54 113.753
R2833 a_27762_11446.t21 a_27762_11446.t12 113.753
R2834 a_27762_11446.t21 a_27762_11446.t24 113.753
R2835 a_27762_11446.t11 a_27762_11446.t14 113.753
R2836 a_27762_11446.t11 a_27762_11446.t27 113.753
R2837 a_27762_11446.t11 a_27762_11446.t40 113.753
R2838 a_27762_11446.t11 a_27762_11446.t56 113.753
R2839 a_27762_11446.t21 a_27762_11446.t49 113.753
R2840 a_27762_11446.t21 a_27762_11446.t4 113.753
R2841 a_27762_11446.t21 a_27762_11446.t19 113.753
R2842 a_27762_11446.t21 a_27762_11446.t34 113.753
R2843 a_27762_11446.t11 a_27762_11446.t48 113.753
R2844 a_27762_11446.t11 a_27762_11446.t2 113.753
R2845 a_27762_11446.t11 a_27762_11446.t18 113.753
R2846 a_27762_11446.t11 a_27762_11446.t33 113.753
R2847 a_27762_11446.n0 a_27762_11446.t11 88.886
R2848 a_27762_11446.n0 a_27762_11446.t1 81.996
R2849 a_27762_11446.t0 a_27762_11446.n0 59.267
R2850 a_27762_11446.t11 a_27762_11446.t21 23.892
R2851 a_28994_11501.n0 a_28994_11501.n6 75.709
R2852 a_28994_11501.n4 a_28994_11501.n5 75.708
R2853 a_28994_11501.n1 a_28994_11501.n2 75.707
R2854 a_28994_11501.n2 a_28994_11501.n3 75.707
R2855 a_28994_11501.n3 a_28994_11501.n4 75.707
R2856 a_28994_11501.n0 a_28994_11501.n1 75.706
R2857 a_28994_11501.n0 a_28994_11501.t5 17.401
R2858 a_28994_11501.n4 a_28994_11501.t3 17.401
R2859 a_28994_11501.n3 a_28994_11501.t7 17.401
R2860 a_28994_11501.n2 a_28994_11501.t4 17.401
R2861 a_28994_11501.n1 a_28994_11501.t2 17.401
R2862 a_28994_11501.n5 a_28994_11501.t6 17.4
R2863 a_28994_11501.n5 a_28994_11501.t13 17.4
R2864 a_28994_11501.n4 a_28994_11501.t11 17.4
R2865 a_28994_11501.n3 a_28994_11501.t12 17.4
R2866 a_28994_11501.n2 a_28994_11501.t10 17.4
R2867 a_28994_11501.n1 a_28994_11501.t9 17.4
R2868 a_28994_11501.n6 a_28994_11501.t8 17.4
R2869 a_28994_11501.n6 a_28994_11501.t1 17.4
R2870 a_28994_11501.t0 a_28994_11501.n0 17.4
R2871 a_29252_11501.n0 a_29252_11501.n6 75.709
R2872 a_29252_11501.n4 a_29252_11501.n5 75.708
R2873 a_29252_11501.n1 a_29252_11501.n2 75.707
R2874 a_29252_11501.n2 a_29252_11501.n3 75.707
R2875 a_29252_11501.n3 a_29252_11501.n4 75.707
R2876 a_29252_11501.n0 a_29252_11501.n1 75.706
R2877 a_29252_11501.n0 a_29252_11501.t1 17.401
R2878 a_29252_11501.n4 a_29252_11501.t3 17.401
R2879 a_29252_11501.n3 a_29252_11501.t5 17.401
R2880 a_29252_11501.n2 a_29252_11501.t4 17.401
R2881 a_29252_11501.n1 a_29252_11501.t6 17.401
R2882 a_29252_11501.n5 a_29252_11501.t0 17.4
R2883 a_29252_11501.n5 a_29252_11501.t7 17.4
R2884 a_29252_11501.n4 a_29252_11501.t10 17.4
R2885 a_29252_11501.n3 a_29252_11501.t8 17.4
R2886 a_29252_11501.n2 a_29252_11501.t11 17.4
R2887 a_29252_11501.n1 a_29252_11501.t9 17.4
R2888 a_29252_11501.n6 a_29252_11501.t2 17.4
R2889 a_29252_11501.n6 a_29252_11501.t13 17.4
R2890 a_29252_11501.t12 a_29252_11501.n0 17.4
R2891 a_49932_4124.t2 a_49932_4124.n0 13.614
R2892 a_49932_4124.n0 a_49932_4124.t3 8.097
R2893 a_49932_4124.n0 a_49932_4124.n1 3.595
R2894 a_49932_4124.n1 a_49932_4124.t1 33.597
R2895 a_49932_4124.n1 a_49932_4124.t0 1.976
R2896 a_65088_25280.n0 a_65088_25280.t5 203.459
R2897 a_65088_25280.n1 a_65088_25280.t3 187.847
R2898 a_65088_25280.n1 a_65088_25280.t2 164.979
R2899 a_65088_25280.n0 a_65088_25280.t4 149.105
R2900 a_65088_25280.n3 a_65088_25280.t1 143.732
R2901 a_65088_25280.n2 a_65088_25280.n1 76
R2902 a_65088_25280.t0 a_65088_25280.n3 73.482
R2903 a_65088_25280.n3 a_65088_25280.n2 50.925
R2904 a_65088_25280.n2 a_65088_25280.n0 41.551
R2905 a_65343_25280.n1 a_65343_25280.n0 163.71
R2906 a_65343_25280.t0 a_65343_25280.n1 82.083
R2907 a_65343_25280.n0 a_65343_25280.t3 63.333
R2908 a_65343_25280.n1 a_65343_25280.t2 63.321
R2909 a_65343_25280.n0 a_65343_25280.t1 29.726
R2910 a_65438_25280.n1 a_65438_25280.t4 332.579
R2911 a_65438_25280.n1 a_65438_25280.t5 168.699
R2912 a_65438_25280.n2 a_65438_25280.n1 104.381
R2913 a_65438_25280.n2 a_65438_25280.n0 101.869
R2914 a_65438_25280.t0 a_65438_25280.n3 96.154
R2915 a_65438_25280.n3 a_65438_25280.n2 92.648
R2916 a_65438_25280.n3 a_65438_25280.t2 65.666
R2917 a_65438_25280.n0 a_65438_25280.t3 65
R2918 a_65438_25280.n0 a_65438_25280.t1 45
R2919 a_66346_26048.t0 a_66346_26048.t1 87.142
R2920 a_26331_5596.n0 a_26331_5596.n1 75.71
R2921 a_26331_5596.n4 a_26331_5596.n5 75.708
R2922 a_26331_5596.n2 a_26331_5596.n3 75.707
R2923 a_26331_5596.n3 a_26331_5596.n4 75.707
R2924 a_26331_5596.n1 a_26331_5596.n6 75.707
R2925 a_26331_5596.n0 a_26331_5596.n2 75.706
R2926 a_26331_5596.t6 a_26331_5596.n0 17.401
R2927 a_26331_5596.n4 a_26331_5596.t0 17.401
R2928 a_26331_5596.n3 a_26331_5596.t5 17.401
R2929 a_26331_5596.n2 a_26331_5596.t1 17.401
R2930 a_26331_5596.n1 a_26331_5596.t4 17.401
R2931 a_26331_5596.n5 a_26331_5596.t3 17.4
R2932 a_26331_5596.n5 a_26331_5596.t11 17.4
R2933 a_26331_5596.n4 a_26331_5596.t12 17.4
R2934 a_26331_5596.n3 a_26331_5596.t8 17.4
R2935 a_26331_5596.n2 a_26331_5596.t13 17.4
R2936 a_26331_5596.n1 a_26331_5596.t7 17.4
R2937 a_26331_5596.n6 a_26331_5596.t2 17.4
R2938 a_26331_5596.n6 a_26331_5596.t10 17.4
R2939 a_26331_5596.n0 a_26331_5596.t9 17.4
R2940 a_65656_25522.n1 a_65656_25522.t5 350.253
R2941 a_65656_25522.n1 a_65656_25522.t4 189.586
R2942 a_65656_25522.n2 a_65656_25522.n1 97.205
R2943 a_65656_25522.n3 a_65656_25522.t3 89.119
R2944 a_65656_25522.n2 a_65656_25522.n0 79.305
R2945 a_65656_25522.n3 a_65656_25522.n2 66.705
R2946 a_65656_25522.n0 a_65656_25522.t2 63.333
R2947 a_65656_25522.t1 a_65656_25522.n3 41.041
R2948 a_65656_25522.n0 a_65656_25522.t0 31.979
R2949 a_44752_16348.t2 a_44752_16348.n2 349.137
R2950 a_44752_16348.n1 a_44752_16348.t4 197.553
R2951 a_44752_16348.n0 a_44752_16348.t1 178.539
R2952 a_44752_16348.n0 a_44752_16348.t3 122.603
R2953 a_44752_16348.n1 a_44752_16348.t0 114.713
R2954 a_44752_16348.n2 a_44752_16348.n0 95.215
R2955 a_44752_16348.n2 a_44752_16348.n1 26.034
R2956 a_51138_19904.t0 a_51138_19904.n0 171.568
R2957 a_51138_19904.n0 a_51138_19904.t2 171.564
R2958 a_51138_19904.n0 a_51138_19904.t1 171.52
R2959 a_25557_17217.n4 a_25557_17217.n5 75.437
R2960 a_25557_17217.n0 a_25557_17217.n1 75.436
R2961 a_25557_17217.n1 a_25557_17217.n2 75.436
R2962 a_25557_17217.n2 a_25557_17217.n3 75.436
R2963 a_25557_17217.n3 a_25557_17217.n4 75.436
R2964 a_25557_17217.n6 a_25557_17217.n0 75.436
R2965 a_25557_17217.n4 a_25557_17217.t0 17.401
R2966 a_25557_17217.n3 a_25557_17217.t13 17.401
R2967 a_25557_17217.n2 a_25557_17217.t11 17.401
R2968 a_25557_17217.n1 a_25557_17217.t9 17.401
R2969 a_25557_17217.n0 a_25557_17217.t10 17.401
R2970 a_25557_17217.n5 a_25557_17217.t12 17.4
R2971 a_25557_17217.n5 a_25557_17217.t1 17.4
R2972 a_25557_17217.n4 a_25557_17217.t5 17.4
R2973 a_25557_17217.n3 a_25557_17217.t2 17.4
R2974 a_25557_17217.n2 a_25557_17217.t6 17.4
R2975 a_25557_17217.n1 a_25557_17217.t4 17.4
R2976 a_25557_17217.n0 a_25557_17217.t3 17.4
R2977 a_25557_17217.n6 a_25557_17217.t8 17.4
R2978 a_25557_17217.t7 a_25557_17217.n6 17.4
R2979 a_27962_11501.n6 a_27962_11501.n4 75.711
R2980 a_27962_11501.n1 a_27962_11501.n0 75.707
R2981 a_27962_11501.n2 a_27962_11501.n1 75.707
R2982 a_27962_11501.n3 a_27962_11501.n2 75.707
R2983 a_27962_11501.n4 a_27962_11501.n3 75.707
R2984 a_27962_11501.n0 a_27962_11501.n5 75.707
R2985 a_27962_11501.n4 a_27962_11501.t13 17.401
R2986 a_27962_11501.n3 a_27962_11501.t10 17.401
R2987 a_27962_11501.n2 a_27962_11501.t8 17.401
R2988 a_27962_11501.n1 a_27962_11501.t9 17.401
R2989 a_27962_11501.n0 a_27962_11501.t12 17.401
R2990 a_27962_11501.n4 a_27962_11501.t2 17.4
R2991 a_27962_11501.n3 a_27962_11501.t0 17.4
R2992 a_27962_11501.n2 a_27962_11501.t3 17.4
R2993 a_27962_11501.n1 a_27962_11501.t1 17.4
R2994 a_27962_11501.n0 a_27962_11501.t4 17.4
R2995 a_27962_11501.n5 a_27962_11501.t11 17.4
R2996 a_27962_11501.n5 a_27962_11501.t5 17.4
R2997 a_27962_11501.n6 a_27962_11501.t7 17.4
R2998 a_27962_11501.t6 a_27962_11501.n6 17.4
R2999 a_14832_12082.n1 a_14832_12082.t3 434.515
R3000 a_14832_12082.n0 a_14832_12082.t2 217.163
R3001 a_14832_12082.t1 a_14832_12082.n1 52.152
R3002 a_14832_12082.n0 a_14832_12082.t0 3.106
R3003 a_14832_12082.n1 a_14832_12082.n0 0.908
R3004 CLK_BY_4_IPH_BAR.n1 CLK_BY_4_IPH_BAR.t3 449.587
R3005 CLK_BY_4_IPH_BAR.n1 CLK_BY_4_IPH_BAR.t0 402.739
R3006 CLK_BY_4_IPH_BAR.n0 CLK_BY_4_IPH_BAR.t1 270.989
R3007 CLK_BY_4_IPH_BAR.n0 CLK_BY_4_IPH_BAR.t2 227.612
R3008 CLK_BY_4_IPH_BAR.n2 CLK_BY_4_IPH_BAR.n0 199.119
R3009 CLK_BY_4_IPH_BAR CLK_BY_4_IPH_BAR.n2 155.826
R3010 CLK_BY_4_IPH_BAR.n2 CLK_BY_4_IPH_BAR.n1 38.57
R3011 zz.n1 zz.t0 23.439
R3012 zz.n1 zz.n0 159.637
R3013 zz.n2 zz.n1 5.413
R3014 zz.n3 zz.n4 1.634
R3015 zz.n3 zz.n2 0.549
R3016 zz.n4 zz.t1 19.8
R3017 zz.n4 zz.t2 19.8
R3018 zz zz.n3 5.731
R3019 zz.n2 zz.t3 27.204
R3020 a_64922_25280.n3 a_64922_25280.t5 530.008
R3021 a_64922_25280.n2 a_64922_25280.t2 334.888
R3022 a_64922_25280.n7 a_64922_25280.t7 255.459
R3023 a_64922_25280.n5 a_64922_25280.t4 224.611
R3024 a_64922_25280.n2 a_64922_25280.t6 196.882
R3025 a_64922_25280.n3 a_64922_25280.t3 141.921
R3026 a_64922_25280.t0 a_64922_25280.n8 126.03
R3027 a_64922_25280.n0 a_64922_25280.t1 99.672
R3028 a_64922_25280.n4 a_64922_25280.n3 92.562
R3029 a_64922_25280.n4 a_64922_25280.n2 44.57
R3030 a_64922_25280.n0 a_64922_25280.n4 38.638
R3031 a_64922_25280.n1 a_64922_25280.n6 15
R3032 a_64922_25280.n8 a_64922_25280.n7 15
R3033 a_64922_25280.n1 a_64922_25280.n5 13.653
R3034 a_64922_25280.n8 a_64922_25280.n1 3.182
R3035 a_64922_25280.n1 a_64922_25280.n0 2.692
R3036 a_66003_25280.n1 a_66003_25280.t5 366.855
R3037 a_66003_25280.n1 a_66003_25280.t4 174.055
R3038 a_66003_25280.n2 a_66003_25280.n0 117.298
R3039 a_66003_25280.n2 a_66003_25280.n1 77.111
R3040 a_66003_25280.n0 a_66003_25280.t3 70
R3041 a_66003_25280.t1 a_66003_25280.n3 68.011
R3042 a_66003_25280.n3 a_66003_25280.t2 63.321
R3043 a_66003_25280.n0 a_66003_25280.t0 61.666
R3044 a_66003_25280.n3 a_66003_25280.n2 57.017
R3045 a_56334_19906.t0 a_56334_19906.t1 343.04
R3046 a_26073_5596.n0 a_26073_5596.n1 75.71
R3047 a_26073_5596.n4 a_26073_5596.n5 75.708
R3048 a_26073_5596.n2 a_26073_5596.n3 75.707
R3049 a_26073_5596.n3 a_26073_5596.n4 75.707
R3050 a_26073_5596.n1 a_26073_5596.n6 75.707
R3051 a_26073_5596.n0 a_26073_5596.n2 75.706
R3052 a_26073_5596.t6 a_26073_5596.n0 17.401
R3053 a_26073_5596.n4 a_26073_5596.t0 17.401
R3054 a_26073_5596.n3 a_26073_5596.t5 17.401
R3055 a_26073_5596.n2 a_26073_5596.t1 17.401
R3056 a_26073_5596.n1 a_26073_5596.t4 17.401
R3057 a_26073_5596.n5 a_26073_5596.t3 17.4
R3058 a_26073_5596.n5 a_26073_5596.t11 17.4
R3059 a_26073_5596.n4 a_26073_5596.t8 17.4
R3060 a_26073_5596.n3 a_26073_5596.t13 17.4
R3061 a_26073_5596.n2 a_26073_5596.t9 17.4
R3062 a_26073_5596.n1 a_26073_5596.t12 17.4
R3063 a_26073_5596.n6 a_26073_5596.t2 17.4
R3064 a_26073_5596.n6 a_26073_5596.t10 17.4
R3065 a_26073_5596.n0 a_26073_5596.t7 17.4
R3066 a_23919_17217.n0 a_23919_17217.n2 75.71
R3067 a_23919_17217.n4 a_23919_17217.n5 75.708
R3068 a_23919_17217.n2 a_23919_17217.n1 75.707
R3069 a_23919_17217.n3 a_23919_17217.n4 75.707
R3070 a_23919_17217.n1 a_23919_17217.n6 75.707
R3071 a_23919_17217.n0 a_23919_17217.n3 75.706
R3072 a_23919_17217.t0 a_23919_17217.n0 17.401
R3073 a_23919_17217.n4 a_23919_17217.t4 17.401
R3074 a_23919_17217.n3 a_23919_17217.t7 17.401
R3075 a_23919_17217.n2 a_23919_17217.t3 17.401
R3076 a_23919_17217.n1 a_23919_17217.t8 17.401
R3077 a_23919_17217.n5 a_23919_17217.t9 17.4
R3078 a_23919_17217.n5 a_23919_17217.t2 17.4
R3079 a_23919_17217.n4 a_23919_17217.t11 17.4
R3080 a_23919_17217.n3 a_23919_17217.t12 17.4
R3081 a_23919_17217.n2 a_23919_17217.t10 17.4
R3082 a_23919_17217.n1 a_23919_17217.t13 17.4
R3083 a_23919_17217.n6 a_23919_17217.t1 17.4
R3084 a_23919_17217.n6 a_23919_17217.t6 17.4
R3085 a_23919_17217.n0 a_23919_17217.t5 17.4
R3086 a_24177_17217.n4 a_24177_17217.n5 75.708
R3087 a_24177_17217.n0 a_24177_17217.n1 75.707
R3088 a_24177_17217.n1 a_24177_17217.n2 75.707
R3089 a_24177_17217.n2 a_24177_17217.n3 75.707
R3090 a_24177_17217.n3 a_24177_17217.n4 75.707
R3091 a_24177_17217.n6 a_24177_17217.n0 75.707
R3092 a_24177_17217.n4 a_24177_17217.t11 17.401
R3093 a_24177_17217.n3 a_24177_17217.t12 17.401
R3094 a_24177_17217.n2 a_24177_17217.t1 17.401
R3095 a_24177_17217.n1 a_24177_17217.t3 17.401
R3096 a_24177_17217.n0 a_24177_17217.t2 17.401
R3097 a_24177_17217.n5 a_24177_17217.t13 17.4
R3098 a_24177_17217.n5 a_24177_17217.t4 17.4
R3099 a_24177_17217.n4 a_24177_17217.t8 17.4
R3100 a_24177_17217.n3 a_24177_17217.t5 17.4
R3101 a_24177_17217.n2 a_24177_17217.t9 17.4
R3102 a_24177_17217.n1 a_24177_17217.t7 17.4
R3103 a_24177_17217.n0 a_24177_17217.t6 17.4
R3104 a_24177_17217.n6 a_24177_17217.t0 17.4
R3105 a_24177_17217.t10 a_24177_17217.n6 17.4
R3106 a_23160_10936.n0 a_23160_10936.t0 391.966
R3107 a_23160_10936.t6 a_23160_10936.n5 93.107
R3108 a_23160_10936.n1 a_23160_10936.n0 75.707
R3109 a_23160_10936.n5 a_23160_10936.n4 75.707
R3110 a_23160_10936.n4 a_23160_10936.n3 75.707
R3111 a_23160_10936.n3 a_23160_10936.n2 75.707
R3112 a_23160_10936.n2 a_23160_10936.n1 75.707
R3113 a_23160_10936.n0 a_23160_10936.t7 17.401
R3114 a_23160_10936.n1 a_23160_10936.t3 17.401
R3115 a_23160_10936.n2 a_23160_10936.t1 17.401
R3116 a_23160_10936.n3 a_23160_10936.t4 17.401
R3117 a_23160_10936.n4 a_23160_10936.t2 17.401
R3118 a_23160_10936.n5 a_23160_10936.t5 17.401
R3119 Vso7b.n0 Vso7b.t1 17.996
R3120 Vso7b Vso7b.n1 0.176
R3121 Vso7b.n1 Vso7b.n0 1.272
R3122 Vso7b.n1 Vso7b.n4 7.169
R3123 Vso7b.n4 Vso7b.t3 420.39
R3124 Vso7b.n4 Vso7b.n3 154.461
R3125 Vso7b.n3 Vso7b.t5 293.485
R3126 Vso7b.n3 Vso7b.n2 61
R3127 Vso7b.n2 Vso7b.t2 381.726
R3128 Vso7b.n2 Vso7b.t4 385.214
R3129 Vso7b.n0 Vso7b.t0 132.37
R3130 a_8748_11114.t0 a_8748_11114.t1 53.512
R3131 a_23403_11500.n0 a_23403_11500.n2 75.71
R3132 a_23403_11500.n4 a_23403_11500.n5 75.708
R3133 a_23403_11500.n2 a_23403_11500.n1 75.707
R3134 a_23403_11500.n3 a_23403_11500.n4 75.707
R3135 a_23403_11500.n1 a_23403_11500.n6 75.707
R3136 a_23403_11500.n0 a_23403_11500.n3 75.706
R3137 a_23403_11500.t0 a_23403_11500.n0 17.401
R3138 a_23403_11500.n4 a_23403_11500.t2 17.401
R3139 a_23403_11500.n3 a_23403_11500.t3 17.401
R3140 a_23403_11500.n2 a_23403_11500.t4 17.401
R3141 a_23403_11500.n1 a_23403_11500.t1 17.401
R3142 a_23403_11500.n5 a_23403_11500.t6 17.4
R3143 a_23403_11500.n5 a_23403_11500.t12 17.4
R3144 a_23403_11500.n4 a_23403_11500.t10 17.4
R3145 a_23403_11500.n3 a_23403_11500.t13 17.4
R3146 a_23403_11500.n2 a_23403_11500.t7 17.4
R3147 a_23403_11500.n1 a_23403_11500.t8 17.4
R3148 a_23403_11500.n6 a_23403_11500.t5 17.4
R3149 a_23403_11500.n6 a_23403_11500.t9 17.4
R3150 a_23403_11500.n0 a_23403_11500.t11 17.4
R3151 a_23661_11500.n4 a_23661_11500.n5 75.708
R3152 a_23661_11500.n0 a_23661_11500.n1 75.707
R3153 a_23661_11500.n1 a_23661_11500.n2 75.707
R3154 a_23661_11500.n2 a_23661_11500.n3 75.707
R3155 a_23661_11500.n3 a_23661_11500.n4 75.707
R3156 a_23661_11500.n6 a_23661_11500.n0 75.707
R3157 a_23661_11500.n4 a_23661_11500.t3 17.401
R3158 a_23661_11500.n3 a_23661_11500.t1 17.401
R3159 a_23661_11500.n2 a_23661_11500.t4 17.401
R3160 a_23661_11500.n1 a_23661_11500.t2 17.401
R3161 a_23661_11500.n0 a_23661_11500.t5 17.401
R3162 a_23661_11500.n5 a_23661_11500.t0 17.4
R3163 a_23661_11500.n5 a_23661_11500.t11 17.4
R3164 a_23661_11500.n4 a_23661_11500.t7 17.4
R3165 a_23661_11500.n3 a_23661_11500.t12 17.4
R3166 a_23661_11500.n2 a_23661_11500.t8 17.4
R3167 a_23661_11500.n1 a_23661_11500.t13 17.4
R3168 a_23661_11500.n0 a_23661_11500.t9 17.4
R3169 a_23661_11500.t6 a_23661_11500.n6 17.4
R3170 a_23661_11500.n6 a_23661_11500.t10 17.4
R3171 a_42550_16062.t1 a_42550_16062.n0 14.302
R3172 a_42550_16062.n3 a_42550_16062.t2 17.453
R3173 a_42550_16062.n0 a_42550_16062.n3 1.627
R3174 a_42550_16062.n3 a_42550_16062.t0 17.451
R3175 a_42550_16062.n0 a_42550_16062.n2 0.036
R3176 a_42550_16062.n2 a_42550_16062.t3 14.437
R3177 a_42550_16062.n2 a_42550_16062.n1 65.242
R3178 a_42550_16062.n1 a_42550_16062.t4 142.533
R3179 a_42550_16062.n1 a_42550_16062.t5 142.195
R3180 a_42574_15624.t2 a_42574_15624.n4 17.598
R3181 a_42574_15624.n2 a_42574_15624.n3 1.885
R3182 a_42574_15624.n4 a_42574_15624.n2 1.609
R3183 a_42574_15624.n3 a_42574_15624.t3 18.036
R3184 a_42574_15624.n3 a_42574_15624.t1 17.538
R3185 a_42574_15624.n2 a_42574_15624.t4 14.302
R3186 a_42574_15624.n4 a_42574_15624.n1 43.347
R3187 a_42574_15624.n1 a_42574_15624.n0 891.943
R3188 a_42574_15624.n0 a_42574_15624.t5 5.713
R3189 a_42574_15624.n0 a_42574_15624.t0 5.713
R3190 a_42574_15624.n1 a_42574_15624.t6 533.962
R3191 vbiasr vbiasr.t0 3.733
R3192 a_53308_3580.t0 a_53308_3580.t1 7.204
R3193 a_23403_17217.n0 a_23403_17217.n3 75.71
R3194 a_23403_17217.n4 a_23403_17217.n5 75.708
R3195 a_23403_17217.n2 a_23403_17217.n1 75.707
R3196 a_23403_17217.n3 a_23403_17217.n2 75.707
R3197 a_23403_17217.n1 a_23403_17217.n6 75.707
R3198 a_23403_17217.n0 a_23403_17217.n4 75.706
R3199 a_23403_17217.n0 a_23403_17217.t2 17.401
R3200 a_23403_17217.n4 a_23403_17217.t6 17.401
R3201 a_23403_17217.n3 a_23403_17217.t3 17.401
R3202 a_23403_17217.n2 a_23403_17217.t5 17.401
R3203 a_23403_17217.n1 a_23403_17217.t0 17.401
R3204 a_23403_17217.n5 a_23403_17217.t1 17.4
R3205 a_23403_17217.n5 a_23403_17217.t11 17.4
R3206 a_23403_17217.n4 a_23403_17217.t8 17.4
R3207 a_23403_17217.n3 a_23403_17217.t9 17.4
R3208 a_23403_17217.n2 a_23403_17217.t7 17.4
R3209 a_23403_17217.n1 a_23403_17217.t13 17.4
R3210 a_23403_17217.n6 a_23403_17217.t4 17.4
R3211 a_23403_17217.n6 a_23403_17217.t10 17.4
R3212 a_23403_17217.t12 a_23403_17217.n0 17.4
R3213 a_23661_17217.n4 a_23661_17217.n5 75.708
R3214 a_23661_17217.n0 a_23661_17217.n1 75.707
R3215 a_23661_17217.n1 a_23661_17217.n2 75.707
R3216 a_23661_17217.n2 a_23661_17217.n3 75.707
R3217 a_23661_17217.n3 a_23661_17217.n4 75.707
R3218 a_23661_17217.n6 a_23661_17217.n0 75.707
R3219 a_23661_17217.n4 a_23661_17217.t4 17.401
R3220 a_23661_17217.n3 a_23661_17217.t1 17.401
R3221 a_23661_17217.n2 a_23661_17217.t5 17.401
R3222 a_23661_17217.n1 a_23661_17217.t3 17.401
R3223 a_23661_17217.n0 a_23661_17217.t2 17.401
R3224 a_23661_17217.n5 a_23661_17217.t0 17.4
R3225 a_23661_17217.n5 a_23661_17217.t11 17.4
R3226 a_23661_17217.n4 a_23661_17217.t8 17.4
R3227 a_23661_17217.n3 a_23661_17217.t12 17.4
R3228 a_23661_17217.n2 a_23661_17217.t9 17.4
R3229 a_23661_17217.n1 a_23661_17217.t7 17.4
R3230 a_23661_17217.n0 a_23661_17217.t13 17.4
R3231 a_23661_17217.t6 a_23661_17217.n6 17.4
R3232 a_23661_17217.n6 a_23661_17217.t10 17.4
R3233 a_22887_11500.n4 a_22887_11500.n5 75.437
R3234 a_22887_11500.n0 a_22887_11500.n1 75.436
R3235 a_22887_11500.n1 a_22887_11500.n2 75.436
R3236 a_22887_11500.n2 a_22887_11500.n3 75.436
R3237 a_22887_11500.n3 a_22887_11500.n4 75.436
R3238 a_22887_11500.n6 a_22887_11500.n0 75.436
R3239 a_22887_11500.n4 a_22887_11500.t8 17.401
R3240 a_22887_11500.n3 a_22887_11500.t13 17.401
R3241 a_22887_11500.n2 a_22887_11500.t11 17.401
R3242 a_22887_11500.n1 a_22887_11500.t7 17.401
R3243 a_22887_11500.n0 a_22887_11500.t12 17.401
R3244 a_22887_11500.n5 a_22887_11500.t10 17.4
R3245 a_22887_11500.n5 a_22887_11500.t0 17.4
R3246 a_22887_11500.n4 a_22887_11500.t3 17.4
R3247 a_22887_11500.n3 a_22887_11500.t1 17.4
R3248 a_22887_11500.n2 a_22887_11500.t4 17.4
R3249 a_22887_11500.n1 a_22887_11500.t2 17.4
R3250 a_22887_11500.n0 a_22887_11500.t5 17.4
R3251 a_22887_11500.n6 a_22887_11500.t9 17.4
R3252 a_22887_11500.t6 a_22887_11500.n6 17.4
R3253 a_66742_25280.n0 a_66742_25280.t2 239.038
R3254 a_66742_25280.n0 a_66742_25280.t3 166.738
R3255 a_66742_25280.t0 a_66742_25280.n1 95.895
R3256 a_66742_25280.n1 a_66742_25280.t1 71.217
R3257 a_66742_25280.n1 a_66742_25280.n0 30.051
R3258 a_29510_11501.n4 a_29510_11501.n5 75.708
R3259 a_29510_11501.n0 a_29510_11501.n1 75.707
R3260 a_29510_11501.n1 a_29510_11501.n2 75.707
R3261 a_29510_11501.n2 a_29510_11501.n3 75.707
R3262 a_29510_11501.n3 a_29510_11501.n4 75.707
R3263 a_29510_11501.n6 a_29510_11501.n0 75.707
R3264 a_29510_11501.n4 a_29510_11501.t4 17.401
R3265 a_29510_11501.n3 a_29510_11501.t1 17.401
R3266 a_29510_11501.n2 a_29510_11501.t5 17.401
R3267 a_29510_11501.n1 a_29510_11501.t6 17.401
R3268 a_29510_11501.n0 a_29510_11501.t2 17.401
R3269 a_29510_11501.n5 a_29510_11501.t0 17.4
R3270 a_29510_11501.n5 a_29510_11501.t13 17.4
R3271 a_29510_11501.n4 a_29510_11501.t9 17.4
R3272 a_29510_11501.n3 a_29510_11501.t7 17.4
R3273 a_29510_11501.n2 a_29510_11501.t10 17.4
R3274 a_29510_11501.n1 a_29510_11501.t8 17.4
R3275 a_29510_11501.n0 a_29510_11501.t11 17.4
R3276 a_29510_11501.n6 a_29510_11501.t3 17.4
R3277 a_29510_11501.t12 a_29510_11501.n6 17.4
R3278 a_28438_10874.n0 a_28438_10874.t0 338.927
R3279 a_28438_10874.n2 a_28438_10874.t4 93.107
R3280 a_28438_10874.n5 a_28438_10874.n4 75.71
R3281 a_28438_10874.n1 a_28438_10874.n0 75.708
R3282 a_28438_10874.n3 a_28438_10874.n2 75.707
R3283 a_28438_10874.n4 a_28438_10874.n3 75.707
R3284 a_28438_10874.n5 a_28438_10874.n1 75.706
R3285 a_28438_10874.t6 a_28438_10874.n5 17.401
R3286 a_28438_10874.n0 a_28438_10874.t5 17.401
R3287 a_28438_10874.n1 a_28438_10874.t1 17.401
R3288 a_28438_10874.n4 a_28438_10874.t2 17.401
R3289 a_28438_10874.n3 a_28438_10874.t7 17.401
R3290 a_28438_10874.n2 a_28438_10874.t3 17.401
R3291 a_63407_26048.t0 a_63407_26048.t1 198.571
R3292 a_63573_26048.t0 a_63573_26048.t1 60
R3293 a_14910_6932.n1 a_14910_6932.t3 434.494
R3294 a_14910_6932.n0 a_14910_6932.t2 217.163
R3295 a_14910_6932.t1 a_14910_6932.n1 52.318
R3296 a_14910_6932.n0 a_14910_6932.t0 3.106
R3297 a_14910_6932.n1 a_14910_6932.n0 0.906
R3298 a_28622_16652.n0 a_28622_16652.t7 251.074
R3299 a_28622_16652.n5 a_28622_16652.t2 93.109
R3300 a_28622_16652.n4 a_28622_16652.n3 75.707
R3301 a_28622_16652.n3 a_28622_16652.n2 75.707
R3302 a_28622_16652.n2 a_28622_16652.n1 75.707
R3303 a_28622_16652.n1 a_28622_16652.n0 75.707
R3304 a_28622_16652.n5 a_28622_16652.n4 75.706
R3305 a_28622_16652.t6 a_28622_16652.n5 17.401
R3306 a_28622_16652.n0 a_28622_16652.t3 17.401
R3307 a_28622_16652.n1 a_28622_16652.t0 17.401
R3308 a_28622_16652.n2 a_28622_16652.t4 17.401
R3309 a_28622_16652.n3 a_28622_16652.t1 17.401
R3310 a_28622_16652.n4 a_28622_16652.t5 17.401
R3311 Vso4b.n0 Vso4b.t1 17.996
R3312 Vso4b Vso4b.n0 0.964
R3313 Vso4b Vso4b.n1 11.542
R3314 Vso4b.n1 Vso4b.t4 412.89
R3315 Vso4b.n1 Vso4b.n3 141.062
R3316 Vso4b.n3 Vso4b.t5 289.419
R3317 Vso4b.n3 Vso4b.n2 58.288
R3318 Vso4b.n2 Vso4b.t2 379.015
R3319 Vso4b.n2 Vso4b.t3 387.926
R3320 Vso4b.n0 Vso4b.t0 132.37
R3321 a_8740_12844.t0 a_8740_12844.t1 53.512
R3322 a_4314_11468.t0 a_4314_11468.t1 12.222
R3323 a_4314_11564.t0 a_4314_11564.t1 12.222
R3324 a_4288_11918.t1 a_4288_11918.n0 18.871
R3325 a_4288_11918.n0 a_4288_11918.n1 1.805
R3326 a_4288_11918.n1 a_4288_11918.t0 26.764
R3327 a_4288_11918.n1 a_4288_11918.n2 3.1
R3328 a_4288_11918.n2 a_4288_11918.t4 595.958
R3329 a_4288_11918.n2 a_4288_11918.t3 433.766
R3330 a_4288_11918.n0 a_4288_11918.t2 17.028
R3331 vout.n8 vout.t0 18.112
R3332 vout.n8 vout.n0 0.852
R3333 vout.n0 vout.n1 0.801
R3334 vout.n3 vout.n8 0.268
R3335 vout.n4 vout.t6 18.897
R3336 vout.n5 vout.n4 0.82
R3337 vout.n6 vout.n5 0.798
R3338 vout.n7 vout.n6 0.836
R3339 vout.n3 vout.n7 0.454
R3340 vout.n7 vout.t7 18.028
R3341 vout.n6 vout.t9 18.148
R3342 vout.n5 vout.t8 18.048
R3343 vout.n4 vout.t1 18.271
R3344 vout.n2 vout.n3 2.226
R3345 vout vout.n2 2.153
R3346 vout.n2 vout.t5 6.206
R3347 vout.n1 vout.t4 19.467
R3348 vout.n1 vout.t2 18.087
R3349 vout.n0 vout.t3 18.418
R3350 a_23145_11500.n0 a_23145_11500.n1 75.71
R3351 a_23145_11500.n4 a_23145_11500.n5 75.708
R3352 a_23145_11500.n2 a_23145_11500.n3 75.707
R3353 a_23145_11500.n3 a_23145_11500.n4 75.707
R3354 a_23145_11500.n1 a_23145_11500.n6 75.707
R3355 a_23145_11500.n0 a_23145_11500.n2 75.706
R3356 a_23145_11500.t6 a_23145_11500.n0 17.401
R3357 a_23145_11500.n4 a_23145_11500.t0 17.401
R3358 a_23145_11500.n3 a_23145_11500.t5 17.401
R3359 a_23145_11500.n2 a_23145_11500.t1 17.401
R3360 a_23145_11500.n1 a_23145_11500.t2 17.401
R3361 a_23145_11500.n5 a_23145_11500.t4 17.4
R3362 a_23145_11500.n5 a_23145_11500.t13 17.4
R3363 a_23145_11500.n4 a_23145_11500.t9 17.4
R3364 a_23145_11500.n3 a_23145_11500.t7 17.4
R3365 a_23145_11500.n2 a_23145_11500.t10 17.4
R3366 a_23145_11500.n1 a_23145_11500.t11 17.4
R3367 a_23145_11500.n6 a_23145_11500.t3 17.4
R3368 a_23145_11500.n6 a_23145_11500.t12 17.4
R3369 a_23145_11500.n0 a_23145_11500.t8 17.4
R3370 a_64615_26048.n0 a_64615_26048.t3 239.038
R3371 a_64615_26048.n0 a_64615_26048.t2 166.738
R3372 a_64615_26048.t0 a_64615_26048.n1 95.895
R3373 a_64615_26048.n1 a_64615_26048.t1 71.217
R3374 a_64615_26048.n1 a_64615_26048.n0 30.051
R3375 CLK_BY_2_BAR.n1 CLK_BY_2_BAR.t6 333.651
R3376 CLK_BY_2_BAR.n1 CLK_BY_2_BAR.t9 297.233
R3377 CLK_BY_2_BAR.n4 CLK_BY_2_BAR.t3 294.554
R3378 CLK_BY_2_BAR.n2 CLK_BY_2_BAR.t5 212.079
R3379 CLK_BY_2_BAR.n3 CLK_BY_2_BAR.t2 212.079
R3380 CLK_BY_2_BAR.n4 CLK_BY_2_BAR.t4 211.008
R3381 CLK_BY_2_BAR.n2 CLK_BY_2_BAR.t8 139.779
R3382 CLK_BY_2_BAR.n3 CLK_BY_2_BAR.t7 139.779
R3383 CLK_BY_2_BAR.n5 CLK_BY_2_BAR.t1 102.408
R3384 CLK_BY_2_BAR.n0 CLK_BY_2_BAR.n3 68.902
R3385 CLK_BY_2_BAR.n3 CLK_BY_2_BAR.n2 61.345
R3386 CLK_BY_2_BAR.n0 CLK_BY_2_BAR.t0 54.537
R3387 CLK_BY_2_BAR CLK_BY_2_BAR.n1 49.8
R3388 CLK_BY_2_BAR CLK_BY_2_BAR.n0 19.824
R3389 CLK_BY_2_BAR.n5 CLK_BY_2_BAR.n4 12.821
R3390 CLK_BY_2_BAR.n0 CLK_BY_2_BAR.n5 4.384
R3391 a_26016_10878.n5 a_26016_10878.t7 305.609
R3392 a_26016_10878.n0 a_26016_10878.t5 93.107
R3393 a_26016_10878.n5 a_26016_10878.n4 75.71
R3394 a_26016_10878.n1 a_26016_10878.n0 75.707
R3395 a_26016_10878.n2 a_26016_10878.n1 75.707
R3396 a_26016_10878.n3 a_26016_10878.n2 75.707
R3397 a_26016_10878.n4 a_26016_10878.n3 75.707
R3398 a_26016_10878.t6 a_26016_10878.n5 17.401
R3399 a_26016_10878.n4 a_26016_10878.t2 17.401
R3400 a_26016_10878.n3 a_26016_10878.t0 17.401
R3401 a_26016_10878.n2 a_26016_10878.t3 17.401
R3402 a_26016_10878.n1 a_26016_10878.t1 17.401
R3403 a_26016_10878.n0 a_26016_10878.t4 17.401
R3404 a_22629_17217.n4 a_22629_17217.n5 75.708
R3405 a_22629_17217.n0 a_22629_17217.n1 75.707
R3406 a_22629_17217.n1 a_22629_17217.n2 75.707
R3407 a_22629_17217.n2 a_22629_17217.n3 75.707
R3408 a_22629_17217.n3 a_22629_17217.n4 75.707
R3409 a_22629_17217.n6 a_22629_17217.n0 75.707
R3410 a_22629_17217.n4 a_22629_17217.t11 17.401
R3411 a_22629_17217.n3 a_22629_17217.t8 17.401
R3412 a_22629_17217.n2 a_22629_17217.t12 17.401
R3413 a_22629_17217.n1 a_22629_17217.t10 17.401
R3414 a_22629_17217.n0 a_22629_17217.t9 17.401
R3415 a_22629_17217.n5 a_22629_17217.t7 17.4
R3416 a_22629_17217.n5 a_22629_17217.t0 17.4
R3417 a_22629_17217.n4 a_22629_17217.t4 17.4
R3418 a_22629_17217.n3 a_22629_17217.t1 17.4
R3419 a_22629_17217.n2 a_22629_17217.t5 17.4
R3420 a_22629_17217.n1 a_22629_17217.t3 17.4
R3421 a_22629_17217.n0 a_22629_17217.t2 17.4
R3422 a_22629_17217.n6 a_22629_17217.t13 17.4
R3423 a_22629_17217.t6 a_22629_17217.n6 17.4
R3424 a_64725_25280.n1 a_64725_25280.t5 294.554
R3425 a_64725_25280.n1 a_64725_25280.t4 211.008
R3426 a_64725_25280.n2 a_64725_25280.n1 45.038
R3427 a_64725_25280.n3 a_64725_25280.t2 26.595
R3428 a_64725_25280.t3 a_64725_25280.n3 26.595
R3429 a_64725_25280.n0 a_64725_25280.t0 24.923
R3430 a_64725_25280.n0 a_64725_25280.t1 24.923
R3431 a_64725_25280.n2 a_64725_25280.n0 20.146
R3432 a_64725_25280.n3 a_64725_25280.n2 19.575
R3433 a_25815_11500.n6 a_25815_11500.n4 75.711
R3434 a_25815_11500.n1 a_25815_11500.n0 75.707
R3435 a_25815_11500.n2 a_25815_11500.n1 75.707
R3436 a_25815_11500.n3 a_25815_11500.n2 75.707
R3437 a_25815_11500.n4 a_25815_11500.n3 75.707
R3438 a_25815_11500.n0 a_25815_11500.n5 75.707
R3439 a_25815_11500.n4 a_25815_11500.t2 17.401
R3440 a_25815_11500.n3 a_25815_11500.t0 17.401
R3441 a_25815_11500.n2 a_25815_11500.t3 17.401
R3442 a_25815_11500.n1 a_25815_11500.t1 17.401
R3443 a_25815_11500.n0 a_25815_11500.t4 17.401
R3444 a_25815_11500.n4 a_25815_11500.t9 17.4
R3445 a_25815_11500.n3 a_25815_11500.t7 17.4
R3446 a_25815_11500.n2 a_25815_11500.t10 17.4
R3447 a_25815_11500.n1 a_25815_11500.t8 17.4
R3448 a_25815_11500.n0 a_25815_11500.t11 17.4
R3449 a_25815_11500.n5 a_25815_11500.t5 17.4
R3450 a_25815_11500.n5 a_25815_11500.t12 17.4
R3451 a_25815_11500.t6 a_25815_11500.n6 17.4
R3452 a_25815_11500.n6 a_25815_11500.t13 17.4
R3453 a_54448_7822.t1 a_54448_7822.t0 184.89
R3454 a_24410_25128.n1 a_24410_25128.t3 434.509
R3455 a_24410_25128.n0 a_24410_25128.t2 217.163
R3456 a_24410_25128.t1 a_24410_25128.n1 52.459
R3457 a_24410_25128.n0 a_24410_25128.t0 3.106
R3458 a_24410_25128.n1 a_24410_25128.n0 0.899
R3459 a_28220_11501.n6 a_28220_11501.n4 75.44
R3460 a_28220_11501.n1 a_28220_11501.n0 75.436
R3461 a_28220_11501.n2 a_28220_11501.n1 75.436
R3462 a_28220_11501.n3 a_28220_11501.n2 75.436
R3463 a_28220_11501.n4 a_28220_11501.n3 75.436
R3464 a_28220_11501.n0 a_28220_11501.n5 75.436
R3465 a_28220_11501.n4 a_28220_11501.t4 17.401
R3466 a_28220_11501.n3 a_28220_11501.t3 17.401
R3467 a_28220_11501.n2 a_28220_11501.t2 17.401
R3468 a_28220_11501.n1 a_28220_11501.t5 17.401
R3469 a_28220_11501.n0 a_28220_11501.t13 17.401
R3470 a_28220_11501.n4 a_28220_11501.t8 17.4
R3471 a_28220_11501.n3 a_28220_11501.t6 17.4
R3472 a_28220_11501.n2 a_28220_11501.t9 17.4
R3473 a_28220_11501.n1 a_28220_11501.t7 17.4
R3474 a_28220_11501.n0 a_28220_11501.t10 17.4
R3475 a_28220_11501.n5 a_28220_11501.t1 17.4
R3476 a_28220_11501.n5 a_28220_11501.t11 17.4
R3477 a_28220_11501.n6 a_28220_11501.t0 17.4
R3478 a_28220_11501.t12 a_28220_11501.n6 17.4
R3479 a_28478_11501.n0 a_28478_11501.n1 75.71
R3480 a_28478_11501.n4 a_28478_11501.n5 75.708
R3481 a_28478_11501.n2 a_28478_11501.n3 75.707
R3482 a_28478_11501.n3 a_28478_11501.n4 75.707
R3483 a_28478_11501.n1 a_28478_11501.n6 75.707
R3484 a_28478_11501.n0 a_28478_11501.n2 75.706
R3485 a_28478_11501.n0 a_28478_11501.t5 17.401
R3486 a_28478_11501.n4 a_28478_11501.t0 17.401
R3487 a_28478_11501.n3 a_28478_11501.t13 17.401
R3488 a_28478_11501.n2 a_28478_11501.t3 17.401
R3489 a_28478_11501.n1 a_28478_11501.t2 17.401
R3490 a_28478_11501.n5 a_28478_11501.t4 17.4
R3491 a_28478_11501.n5 a_28478_11501.t10 17.4
R3492 a_28478_11501.n4 a_28478_11501.t6 17.4
R3493 a_28478_11501.n3 a_28478_11501.t11 17.4
R3494 a_28478_11501.n2 a_28478_11501.t7 17.4
R3495 a_28478_11501.n1 a_28478_11501.t8 17.4
R3496 a_28478_11501.n6 a_28478_11501.t1 17.4
R3497 a_28478_11501.n6 a_28478_11501.t9 17.4
R3498 a_28478_11501.t12 a_28478_11501.n0 17.4
R3499 a_23308_802.n1 a_23308_802.t2 434.515
R3500 a_23308_802.n0 a_23308_802.t3 217.163
R3501 a_23308_802.t1 a_23308_802.n1 52.152
R3502 a_23308_802.n0 a_23308_802.t0 3.106
R3503 a_23308_802.n1 a_23308_802.n0 0.908
R3504 a_26110_16652.n0 a_26110_16652.t7 277.494
R3505 a_26110_16652.t6 a_26110_16652.n5 93.107
R3506 a_26110_16652.n5 a_26110_16652.n4 75.707
R3507 a_26110_16652.n4 a_26110_16652.n3 75.707
R3508 a_26110_16652.n3 a_26110_16652.n2 75.707
R3509 a_26110_16652.n2 a_26110_16652.n1 75.707
R3510 a_26110_16652.n1 a_26110_16652.n0 75.707
R3511 a_26110_16652.n0 a_26110_16652.t0 17.401
R3512 a_26110_16652.n1 a_26110_16652.t4 17.401
R3513 a_26110_16652.n2 a_26110_16652.t1 17.401
R3514 a_26110_16652.n3 a_26110_16652.t5 17.401
R3515 a_26110_16652.n4 a_26110_16652.t3 17.401
R3516 a_26110_16652.n5 a_26110_16652.t2 17.401
R3517 a_8744_9386.t0 a_8744_9386.t1 53.512
R3518 a_4226_12188.t1 a_4226_12188.n0 18.871
R3519 a_4226_12188.n1 a_4226_12188.n2 3.215
R3520 a_4226_12188.n1 a_4226_12188.t0 26.765
R3521 a_4226_12188.n0 a_4226_12188.n1 1.805
R3522 a_4226_12188.n2 a_4226_12188.t3 434.881
R3523 a_4226_12188.n2 a_4226_12188.t4 598.238
R3524 a_4226_12188.n0 a_4226_12188.t2 17.028
R3525 a_32948_24994.n1 a_32948_24994.t3 434.487
R3526 a_32948_24994.n0 a_32948_24994.t2 217.163
R3527 a_32948_24994.t1 a_32948_24994.n1 52.153
R3528 a_32948_24994.n0 a_32948_24994.t0 3.106
R3529 a_32948_24994.n1 a_32948_24994.n0 0.887
R3530 a_28790_25040.n1 a_28790_25040.t3 434.517
R3531 a_28790_25040.n0 a_28790_25040.t2 217.163
R3532 a_28790_25040.t1 a_28790_25040.n1 52.317
R3533 a_28790_25040.n0 a_28790_25040.t0 3.106
R3534 a_28790_25040.n1 a_28790_25040.n0 0.907
R3535 Vso2b.n0 Vso2b.t1 17.996
R3536 Vso2b Vso2b.n0 0.352
R3537 Vso2b Vso2b.n1 4.36
R3538 Vso2b.n1 Vso2b.t4 414.561
R3539 Vso2b.n1 Vso2b.n2 126.708
R3540 Vso2b.n2 Vso2b.n3 57.715
R3541 Vso2b.n3 Vso2b.t2 372.915
R3542 Vso2b.n3 Vso2b.t3 376.403
R3543 Vso2b.n2 Vso2b.t5 283.319
R3544 Vso2b.n0 Vso2b.t0 132.37
R3545 a_66731_26048.n0 a_66731_26048.t2 239.038
R3546 a_66731_26048.n0 a_66731_26048.t3 166.738
R3547 a_66731_26048.t1 a_66731_26048.n1 95.895
R3548 a_66731_26048.n1 a_66731_26048.t0 71.217
R3549 a_66731_26048.n1 a_66731_26048.n0 30.051
R3550 a_51334_14126.t1 a_51334_14126.n0 14.302
R3551 a_51334_14126.n0 a_51334_14126.n7 4.438
R3552 a_51334_14126.n7 a_51334_14126.t3 17.451
R3553 a_51334_14126.n7 a_51334_14126.t0 17.452
R3554 a_51334_14126.n0 a_51334_14126.n1 3.405
R3555 a_51334_14126.n1 a_51334_14126.n5 61.168
R3556 a_51334_14126.n6 a_51334_14126.t5 48.21
R3557 a_51334_14126.n6 a_51334_14126.t7 127.084
R3558 a_51334_14126.n5 a_51334_14126.n6 1.418
R3559 a_51334_14126.n5 a_51334_14126.n3 31.793
R3560 a_51334_14126.n4 a_51334_14126.t8 48.21
R3561 a_51334_14126.n4 a_51334_14126.t4 127.084
R3562 a_51334_14126.n3 a_51334_14126.n4 1.418
R3563 a_51334_14126.n2 a_51334_14126.t9 48.21
R3564 a_51334_14126.n2 a_51334_14126.t6 127.084
R3565 a_51334_14126.n3 a_51334_14126.n2 35.06
R3566 a_51334_14126.n1 a_51334_14126.t2 14.331
R3567 z.n0 z.n1 463.355
R3568 z z.n0 20.186
R3569 z.n0 z.t7 9.051
R3570 z.n0 z.t4 8.766
R3571 z.n0 z.t6 8.705
R3572 z.n0 z.t5 8.7
R3573 z.n0 z.t3 8.7
R3574 z.n0 z.t2 8.7
R3575 z.n1 z.t1 5.713
R3576 z.n1 z.t0 5.713
R3577 a_65992_26048.n1 a_65992_26048.t5 366.855
R3578 a_65992_26048.n1 a_65992_26048.t4 174.055
R3579 a_65992_26048.n2 a_65992_26048.n0 117.298
R3580 a_65992_26048.n2 a_65992_26048.n1 77.111
R3581 a_65992_26048.n0 a_65992_26048.t0 70
R3582 a_65992_26048.t1 a_65992_26048.n3 68.011
R3583 a_65992_26048.n3 a_65992_26048.t2 63.321
R3584 a_65992_26048.n0 a_65992_26048.t3 61.666
R3585 a_65992_26048.n3 a_65992_26048.n2 57.017
R3586 Vso6b.n0 Vso6b.t1 17.996
R3587 Vso6b.n1 Vso6b.n0 0.302
R3588 Vso6b Vso6b.n1 0.335
R3589 Vso6b.n1 Vso6b.n2 2.221
R3590 Vso6b.n2 Vso6b.t3 414.027
R3591 Vso6b.n2 Vso6b.n4 136.535
R3592 Vso6b.n4 Vso6b.t4 292.807
R3593 Vso6b.n4 Vso6b.n3 59.644
R3594 Vso6b.n3 Vso6b.t5 379.693
R3595 Vso6b.n3 Vso6b.t2 387.248
R3596 Vso6b.n0 Vso6b.t0 132.37
R3597 a_4226_11804.t0 a_4226_11804.n0 17.028
R3598 a_4226_11804.n0 a_4226_11804.t1 18.871
R3599 a_4226_11804.n0 a_4226_11804.n2 1.812
R3600 a_4226_11804.n1 a_4226_11804.t4 435.371
R3601 a_4226_11804.n2 a_4226_11804.n1 9.162
R3602 a_4226_11804.n1 a_4226_11804.t3 594.041
R3603 a_4226_11804.n2 a_4226_11804.t2 26.805
R3604 a_51532_4150.n0 a_51532_4150.n1 1.438
R3605 a_51532_4150.n1 a_51532_4150.n2 1.94
R3606 a_51532_4150.n2 a_51532_4150.n4 5.632
R3607 a_51532_4150.n4 a_51532_4150.t4 14.994
R3608 a_51532_4150.n4 a_51532_4150.t6 3.653
R3609 a_51532_4150.n3 a_51532_4150.t0 19.231
R3610 a_51532_4150.n2 a_51532_4150.n3 0.07
R3611 a_51532_4150.n3 a_51532_4150.t5 13.856
R3612 a_51532_4150.n1 a_51532_4150.t1 14.151
R3613 a_51532_4150.n0 a_51532_4150.t2 17.234
R3614 a_51532_4150.t3 a_51532_4150.n0 7.827
R3615 a_64911_26048.n3 a_64911_26048.t6 530.008
R3616 a_64911_26048.n2 a_64911_26048.t5 334.888
R3617 a_64911_26048.n7 a_64911_26048.t2 255.459
R3618 a_64911_26048.n5 a_64911_26048.t3 224.611
R3619 a_64911_26048.n2 a_64911_26048.t4 196.882
R3620 a_64911_26048.n3 a_64911_26048.t7 141.921
R3621 a_64911_26048.t1 a_64911_26048.n8 126.03
R3622 a_64911_26048.n0 a_64911_26048.t0 99.672
R3623 a_64911_26048.n4 a_64911_26048.n3 92.562
R3624 a_64911_26048.n4 a_64911_26048.n2 44.57
R3625 a_64911_26048.n0 a_64911_26048.n4 38.638
R3626 a_64911_26048.n1 a_64911_26048.n6 15
R3627 a_64911_26048.n8 a_64911_26048.n7 15
R3628 a_64911_26048.n1 a_64911_26048.n5 13.653
R3629 a_64911_26048.n8 a_64911_26048.n1 3.182
R3630 a_64911_26048.n1 a_64911_26048.n0 2.692
R3631 a_50032_16080.t1 a_50032_16080.t0 414.247
R3632 a_50262_14152.n0 a_50262_14152.t3 14.474
R3633 a_50262_14152.t0 a_50262_14152.n0 14.302
R3634 a_50262_14152.n0 a_50262_14152.n2 0.512
R3635 a_50262_14152.n2 a_50262_14152.n7 1450.42
R3636 a_50262_14152.n7 a_50262_14152.n6 109.291
R3637 a_50262_14152.n6 a_50262_14152.t9 153.199
R3638 a_50262_14152.n6 a_50262_14152.t6 8.703
R3639 a_50262_14152.n3 a_50262_14152.n4 0.003
R3640 a_50262_14152.n7 a_50262_14152.n3 67.916
R3641 a_50262_14152.n3 a_50262_14152.n5 153.01
R3642 a_50262_14152.n5 a_50262_14152.t5 8.7
R3643 a_50262_14152.n5 a_50262_14152.t7 8.7
R3644 a_50262_14152.n4 a_50262_14152.t8 8.7
R3645 a_50262_14152.n4 a_50262_14152.t4 8.7
R3646 a_50262_14152.n1 a_50262_14152.t2 17.453
R3647 a_50262_14152.n2 a_50262_14152.n1 1.115
R3648 a_50262_14152.n1 a_50262_14152.t1 17.451
R3649 a_50511_16072.n0 a_50511_16072.n1 524.893
R3650 a_50511_16072.n0 a_50511_16072.t8 256.935
R3651 a_50511_16072.n0 a_50511_16072.t1 9.092
R3652 a_50511_16072.t5 a_50511_16072.n0 8.763
R3653 a_50511_16072.n0 a_50511_16072.t0 8.705
R3654 a_50511_16072.n0 a_50511_16072.t2 8.7
R3655 a_50511_16072.n0 a_50511_16072.t3 8.7
R3656 a_50511_16072.n0 a_50511_16072.t4 8.7
R3657 a_50511_16072.n1 a_50511_16072.t6 5.844
R3658 a_50511_16072.n1 a_50511_16072.t7 5.744
R3659 a_50511_16072.t8 a_50511_16072.t9 1.22
R3660 a_62961_26048.n0 a_62961_26048.t5 203.459
R3661 a_62961_26048.n1 a_62961_26048.t4 187.847
R3662 a_62961_26048.n1 a_62961_26048.t3 164.979
R3663 a_62961_26048.n0 a_62961_26048.t2 149.105
R3664 a_62961_26048.n3 a_62961_26048.t0 143.732
R3665 a_62961_26048.n2 a_62961_26048.n1 76
R3666 a_62961_26048.t1 a_62961_26048.n3 73.482
R3667 a_62961_26048.n3 a_62961_26048.n2 50.925
R3668 a_62961_26048.n2 a_62961_26048.n0 41.551
R3669 a_63876_26048.n1 a_63876_26048.t5 366.855
R3670 a_63876_26048.n1 a_63876_26048.t4 174.055
R3671 a_63876_26048.n2 a_63876_26048.n0 117.298
R3672 a_63876_26048.n2 a_63876_26048.n1 77.111
R3673 a_63876_26048.n0 a_63876_26048.t3 70
R3674 a_63876_26048.t1 a_63876_26048.n3 68.011
R3675 a_63876_26048.n3 a_63876_26048.t2 63.321
R3676 a_63876_26048.n0 a_63876_26048.t0 61.666
R3677 a_63876_26048.n3 a_63876_26048.n2 57.017
R3678 a_64038_26414.t0 a_64038_26414.t1 126.642
R3679 a_65534_25280.t1 a_65534_25280.t0 198.571
R3680 a_38070_8852.n1 a_38070_8852.t3 434.515
R3681 a_38070_8852.n0 a_38070_8852.t2 217.163
R3682 a_38070_8852.t1 a_38070_8852.n1 52.152
R3683 a_38070_8852.n0 a_38070_8852.t0 3.106
R3684 a_38070_8852.n1 a_38070_8852.n0 0.908
R3685 a_52052_20224.t0 a_52052_20224.t1 343.213
R3686 a_64230_26048.t0 a_64230_26048.t1 87.142
R3687 a_30384_802.n1 a_30384_802.t3 434.478
R3688 a_30384_802.n0 a_30384_802.t2 217.163
R3689 a_30384_802.t1 a_30384_802.n1 52.152
R3690 a_30384_802.n0 a_30384_802.t0 3.106
R3691 a_30384_802.n1 a_30384_802.n0 0.885
R3692 a_4226_11996.t0 a_4226_11996.n0 17.028
R3693 a_4226_11996.n0 a_4226_11996.t2 18.871
R3694 a_4226_11996.n0 a_4226_11996.n1 1.792
R3695 a_4226_11996.n1 a_4226_11996.n2 7.674
R3696 a_4226_11996.n2 a_4226_11996.t3 595.107
R3697 a_4226_11996.n2 a_4226_11996.t4 363.465
R3698 a_4226_11996.n1 a_4226_11996.t1 26.804
R3699 a_4314_11948.t0 a_4314_11948.t1 12.222
R3700 a_4314_12044.t0 a_4314_12044.t1 12.222
R3701 a_54410_8156.t0 a_54410_8156.t1 343.123
R3702 a_23178_16644.n0 a_23178_16644.t0 333.308
R3703 a_23178_16644.n3 a_23178_16644.t7 93.107
R3704 a_23178_16644.n5 a_23178_16644.n4 75.71
R3705 a_23178_16644.n4 a_23178_16644.n3 75.707
R3706 a_23178_16644.n2 a_23178_16644.n1 75.707
R3707 a_23178_16644.n1 a_23178_16644.n0 75.707
R3708 a_23178_16644.n5 a_23178_16644.n2 75.706
R3709 a_23178_16644.t6 a_23178_16644.n5 17.401
R3710 a_23178_16644.n0 a_23178_16644.t1 17.401
R3711 a_23178_16644.n1 a_23178_16644.t5 17.401
R3712 a_23178_16644.n2 a_23178_16644.t2 17.401
R3713 a_23178_16644.n4 a_23178_16644.t4 17.401
R3714 a_23178_16644.n3 a_23178_16644.t3 17.401
R3715 a_50128_8156.t0 a_50128_8156.t1 343.296
R3716 a_53308_2992.t0 a_53308_2992.t1 25.776
R3717 a_8736_14034.t0 a_8736_14034.t1 53.512
R3718 a_64051_26022.n3 a_64051_26022.t7 389.181
R3719 a_64051_26022.n0 a_64051_26022.t5 256.987
R3720 a_64051_26022.n2 a_64051_26022.t4 212.079
R3721 a_64051_26022.n3 a_64051_26022.t8 174.888
R3722 a_64051_26022.n0 a_64051_26022.t3 163.801
R3723 a_64051_26022.n6 a_64051_26022.n5 161.578
R3724 a_64051_26022.n1 a_64051_26022.t6 139.779
R3725 a_64051_26022.n1 a_64051_26022.n0 129.263
R3726 a_64051_26022.n4 a_64051_26022.n3 102.015
R3727 a_64051_26022.n6 a_64051_26022.t2 63.321
R3728 a_64051_26022.t0 a_64051_26022.n6 63.321
R3729 a_64051_26022.n4 a_64051_26022.t1 46.071
R3730 a_64051_26022.n5 a_64051_26022.n2 37.442
R3731 a_64051_26022.n5 a_64051_26022.n4 23.54
R3732 a_64051_26022.n2 a_64051_26022.n1 22.639
R3733 a_65077_26048.n0 a_65077_26048.t3 203.459
R3734 a_65077_26048.n1 a_65077_26048.t5 187.847
R3735 a_65077_26048.n1 a_65077_26048.t2 164.979
R3736 a_65077_26048.n0 a_65077_26048.t4 149.105
R3737 a_65077_26048.n3 a_65077_26048.t0 143.732
R3738 a_65077_26048.n2 a_65077_26048.n1 76
R3739 a_65077_26048.t1 a_65077_26048.n3 73.482
R3740 a_65077_26048.n3 a_65077_26048.n2 50.925
R3741 a_65077_26048.n2 a_65077_26048.n0 41.551
R3742 a_66112_25280.t1 a_66112_25280.t0 94.726
R3743 a_46856_21176.t0 a_46856_21176.t1 343.213
R3744 a_51138_21494.t1 a_51138_21494.t0 501.405
R3745 a_65427_26048.n1 a_65427_26048.t5 332.579
R3746 a_65427_26048.n1 a_65427_26048.t4 168.699
R3747 a_65427_26048.n2 a_65427_26048.n1 104.381
R3748 a_65427_26048.n2 a_65427_26048.n0 101.869
R3749 a_65427_26048.t1 a_65427_26048.n3 96.154
R3750 a_65427_26048.n3 a_65427_26048.n2 92.648
R3751 a_65427_26048.n3 a_65427_26048.t2 65.666
R3752 a_65427_26048.n0 a_65427_26048.t0 65
R3753 a_65427_26048.n0 a_65427_26048.t3 45
R3754 a_65645_26290.n1 a_65645_26290.t5 350.253
R3755 a_65645_26290.n1 a_65645_26290.t4 189.586
R3756 a_65645_26290.n2 a_65645_26290.n1 97.205
R3757 a_65645_26290.n3 a_65645_26290.t0 89.119
R3758 a_65645_26290.n2 a_65645_26290.n0 79.305
R3759 a_65645_26290.n3 a_65645_26290.n2 66.705
R3760 a_65645_26290.n0 a_65645_26290.t3 63.333
R3761 a_65645_26290.t2 a_65645_26290.n3 41.041
R3762 a_65645_26290.n0 a_65645_26290.t1 31.979
R3763 vbiasot.t2 vbiasot.n2 17.477
R3764 vbiasot.n2 vbiasot.t0 55.042
R3765 vbiasot.n1 vbiasot.n2 0.422
R3766 vbiasot.n1 vbiasot.t1 9.343
R3767 vbiasot vbiasot.n1 5.752
R3768 vbiasot vbiasot.n0 4.17
R3769 vbiasot.n0 vbiasot.t3 0.898
R3770 vbiasot.n0 vbiasot.t4 0.811
R3771 a_25815_17217.n4 a_25815_17217.n5 75.708
R3772 a_25815_17217.n0 a_25815_17217.n1 75.707
R3773 a_25815_17217.n1 a_25815_17217.n2 75.707
R3774 a_25815_17217.n2 a_25815_17217.n3 75.707
R3775 a_25815_17217.n3 a_25815_17217.n4 75.707
R3776 a_25815_17217.n6 a_25815_17217.n0 75.707
R3777 a_25815_17217.n4 a_25815_17217.t4 17.401
R3778 a_25815_17217.n3 a_25815_17217.t1 17.401
R3779 a_25815_17217.n2 a_25815_17217.t5 17.401
R3780 a_25815_17217.n1 a_25815_17217.t3 17.401
R3781 a_25815_17217.n0 a_25815_17217.t2 17.401
R3782 a_25815_17217.n5 a_25815_17217.t0 17.4
R3783 a_25815_17217.n5 a_25815_17217.t7 17.4
R3784 a_25815_17217.n4 a_25815_17217.t11 17.4
R3785 a_25815_17217.n3 a_25815_17217.t8 17.4
R3786 a_25815_17217.n2 a_25815_17217.t12 17.4
R3787 a_25815_17217.n1 a_25815_17217.t10 17.4
R3788 a_25815_17217.n0 a_25815_17217.t9 17.4
R3789 a_25815_17217.t6 a_25815_17217.n6 17.4
R3790 a_25815_17217.n6 a_25815_17217.t13 17.4
R3791 a_4288_12110.t0 a_4288_12110.n0 18.871
R3792 a_4288_12110.n1 a_4288_12110.t1 26.765
R3793 a_4288_12110.n1 a_4288_12110.n2 5.994
R3794 a_4288_12110.n0 a_4288_12110.n1 1.802
R3795 a_4288_12110.n2 a_4288_12110.t3 596.593
R3796 a_4288_12110.n2 a_4288_12110.t4 434.118
R3797 a_4288_12110.n0 a_4288_12110.t2 17.028
R3798 a_23504_23306.t0 a_23504_23306.t1 343.982
R3799 a_46856_19268.n0 a_46856_19268.t0 2113.41
R3800 a_46856_19268.n0 a_46856_19268.t2 171.607
R3801 a_46856_19268.t1 a_46856_19268.n0 171.607
R3802 a_47968_16078.t1 a_47968_16078.n0 14.331
R3803 a_47968_16078.n0 a_47968_16078.n3 191.874
R3804 a_47968_16078.n3 a_47968_16078.t5 5.713
R3805 a_47968_16078.n3 a_47968_16078.t4 5.713
R3806 a_47968_16078.n1 a_47968_16078.n2 4.438
R3807 a_47968_16078.n0 a_47968_16078.n1 3.405
R3808 a_47968_16078.n2 a_47968_16078.t0 17.451
R3809 a_47968_16078.n2 a_47968_16078.t2 17.452
R3810 a_47968_16078.n1 a_47968_16078.t3 14.302
R3811 bb.n0 bb.t0 14.302
R3812 bb.n2 bb.n1 0.039
R3813 bb.n6 bb.n5 0.039
R3814 bb.n7 bb.n3 0.001
R3815 bb.n3 bb.n6 0.045
R3816 bb.n6 bb.n2 0.001
R3817 bb.n2 bb.n8 0.045
R3818 bb.n8 bb.n4 0.001
R3819 bb.n4 bb.n0 1.58
R3820 bb.n9 bb.n7 1.034
R3821 bb.n11 bb.n9 12.792
R3822 bb.n11 bb.t2 210.384
R3823 bb bb.n11 21.932
R3824 bb.n9 bb.n10 1167.29
R3825 bb.n10 bb.t5 142.104
R3826 bb.n10 bb.t6 141.443
R3827 bb.n5 bb.t4 17.411
R3828 bb.n1 bb.t1 17.411
R3829 bb.n0 bb.t3 14.473
R3830 a_4226_11612.t0 a_4226_11612.n0 17.028
R3831 a_4226_11612.n0 a_4226_11612.t1 18.871
R3832 a_4226_11612.n0 a_4226_11612.n1 1.79
R3833 a_4226_11612.n1 a_4226_11612.n2 6.997
R3834 a_4226_11612.n2 a_4226_11612.t4 363.47
R3835 a_4226_11612.n2 a_4226_11612.t3 595.089
R3836 a_4226_11612.n1 a_4226_11612.t2 26.804
R3837 aa.n0 aa.t1 14.331
R3838 aa.n1 aa.n0 0.395
R3839 aa.n0 aa.n5 2.815
R3840 aa.n5 aa.t0 17.453
R3841 aa.n5 aa.t3 17.451
R3842 aa.n1 aa.t4 14.505
R3843 aa.n2 aa.n1 0.764
R3844 aa.n3 aa.n2 4.269
R3845 aa aa.n3 20.947
R3846 aa.n3 aa.n4 1294.49
R3847 aa.n4 aa.t5 139.796
R3848 aa.n4 aa.t6 143.751
R3849 aa.n2 aa.t2 12.589
R3850 a_4288_11726.t0 a_4288_11726.n0 18.871
R3851 a_4288_11726.n0 a_4288_11726.n1 1.815
R3852 a_4288_11726.n1 a_4288_11726.n2 6.196
R3853 a_4288_11726.n2 a_4288_11726.t4 433.807
R3854 a_4288_11726.n2 a_4288_11726.t3 597.059
R3855 a_4288_11726.n1 a_4288_11726.t1 26.804
R3856 a_4288_11726.n0 a_4288_11726.t2 17.028
R3857 a_66101_26048.t1 a_66101_26048.t0 94.726
R3858 a_65535_26414.t0 a_65535_26414.n0 194.654
R3859 a_65535_26414.n0 a_65535_26414.t2 168.384
R3860 a_65535_26414.n0 a_65535_26414.t1 63.321
R3861 Vso8b.n0 Vso8b.t1 17.996
R3862 Vso8b Vso8b.n0 0.614
R3863 Vso8b Vso8b.n3 18.252
R3864 Vso8b.n3 Vso8b.t2 422.392
R3865 Vso8b.n3 Vso8b.n2 154.194
R3866 Vso8b.n2 Vso8b.t5 294.841
R3867 Vso8b.n2 Vso8b.n1 58.966
R3868 Vso8b.n1 Vso8b.t4 380.37
R3869 Vso8b.n1 Vso8b.t3 386.57
R3870 Vso8b.n0 Vso8b.t0 132.37
R3871 CLK_BY_2 CLK_BY_2.t0 58.863
R3872 CLK_BY_2 CLK_BY_2.t1 50.3
R3873 a_51826_16054.t1 a_51826_16054.t0 445.429
R3874 a_43010_16058.t0 a_43010_16058.n0 14.331
R3875 a_43010_16058.n0 a_43010_16058.n1 0.393
R3876 a_43010_16058.n0 a_43010_16058.n3 2.815
R3877 a_43010_16058.n3 a_43010_16058.t1 17.453
R3878 a_43010_16058.n3 a_43010_16058.t2 17.451
R3879 a_43010_16058.n1 a_43010_16058.n2 73.167
R3880 a_43010_16058.n2 a_43010_16058.t5 143.889
R3881 a_43010_16058.n2 a_43010_16058.t4 140.839
R3882 a_43010_16058.n1 a_43010_16058.t3 14.505
R3883 a_28736_11501.n0 a_28736_11501.n1 75.71
R3884 a_28736_11501.n4 a_28736_11501.n5 75.708
R3885 a_28736_11501.n2 a_28736_11501.n3 75.707
R3886 a_28736_11501.n3 a_28736_11501.n4 75.707
R3887 a_28736_11501.n1 a_28736_11501.n6 75.707
R3888 a_28736_11501.n0 a_28736_11501.n2 75.706
R3889 a_28736_11501.n0 a_28736_11501.t13 17.401
R3890 a_28736_11501.n4 a_28736_11501.t7 17.401
R3891 a_28736_11501.n3 a_28736_11501.t12 17.401
R3892 a_28736_11501.n2 a_28736_11501.t8 17.401
R3893 a_28736_11501.n1 a_28736_11501.t9 17.401
R3894 a_28736_11501.n5 a_28736_11501.t11 17.4
R3895 a_28736_11501.n5 a_28736_11501.t4 17.4
R3896 a_28736_11501.n4 a_28736_11501.t0 17.4
R3897 a_28736_11501.n3 a_28736_11501.t5 17.4
R3898 a_28736_11501.n2 a_28736_11501.t1 17.4
R3899 a_28736_11501.n1 a_28736_11501.t2 17.4
R3900 a_28736_11501.n6 a_28736_11501.t10 17.4
R3901 a_28736_11501.n6 a_28736_11501.t3 17.4
R3902 a_28736_11501.t6 a_28736_11501.n0 17.4
R3903 a_66165_25646.t0 a_66165_25646.t1 126.642
R3904 a_65332_26048.n1 a_65332_26048.n0 163.71
R3905 a_65332_26048.n0 a_65332_26048.t3 82.083
R3906 a_65332_26048.n1 a_65332_26048.t0 63.333
R3907 a_65332_26048.n0 a_65332_26048.t2 63.321
R3908 a_65332_26048.n2 a_65332_26048.t1 26.393
R3909 a_65332_26048.n3 a_65332_26048.n2 14.4
R3910 a_65332_26048.n2 a_65332_26048.n1 3.333
R3911 a_42782_16060.t2 a_42782_16060.n0 14.331
R3912 a_42782_16060.n0 a_42782_16060.n4 34.012
R3913 a_42782_16060.n4 a_42782_16060.n3 703.99
R3914 a_42782_16060.n3 a_42782_16060.t1 5.713
R3915 a_42782_16060.n3 a_42782_16060.t0 5.713
R3916 a_42782_16060.n4 a_42782_16060.t6 422.85
R3917 a_42782_16060.n1 a_42782_16060.n2 4.438
R3918 a_42782_16060.n0 a_42782_16060.n1 3.405
R3919 a_42782_16060.n2 a_42782_16060.t3 17.451
R3920 a_42782_16060.n2 a_42782_16060.t4 17.452
R3921 a_42782_16060.n1 a_42782_16060.t5 14.302
R3922 a_4314_11660.t0 a_4314_11660.t1 12.222
R3923 a_4314_11756.t0 a_4314_11756.t1 12.222
R3924 a_66178_25254.n5 a_66178_25254.t5 389.181
R3925 a_66178_25254.n1 a_66178_25254.t4 256.987
R3926 a_66178_25254.n3 a_66178_25254.t7 212.079
R3927 a_66178_25254.n5 a_66178_25254.t6 174.888
R3928 a_66178_25254.n1 a_66178_25254.t8 163.801
R3929 a_66178_25254.n4 a_66178_25254.n0 161.578
R3930 a_66178_25254.n2 a_66178_25254.t3 139.779
R3931 a_66178_25254.n2 a_66178_25254.n1 129.263
R3932 a_66178_25254.n6 a_66178_25254.n5 102.015
R3933 a_66178_25254.n0 a_66178_25254.t1 63.321
R3934 a_66178_25254.n0 a_66178_25254.t2 63.321
R3935 a_66178_25254.t0 a_66178_25254.n6 46.071
R3936 a_66178_25254.n4 a_66178_25254.n3 37.442
R3937 a_66178_25254.n6 a_66178_25254.n4 23.54
R3938 a_66178_25254.n3 a_66178_25254.n2 22.639
R3939 a_51138_20858.t0 a_51138_20858.t1 343.039
R3940 a_47760_15642.t0 a_47760_15642.n0 19.207
R3941 a_47760_15642.n0 a_47760_15642.n2 1.566
R3942 a_47760_15642.n3 a_47760_15642.t2 18.036
R3943 a_47760_15642.n2 a_47760_15642.n3 0.282
R3944 a_47760_15642.n3 a_47760_15642.t1 17.538
R3945 a_47760_15642.n1 a_47760_15642.t4 5.847
R3946 a_47760_15642.n2 a_47760_15642.n1 240.762
R3947 a_47760_15642.n1 a_47760_15642.t5 5.744
R3948 a_47760_15642.n0 a_47760_15642.t3 14.302
R3949 a_8752_10532.t0 a_8752_10532.t1 53.512
R3950 a_4314_12140.t0 a_4314_12140.t1 12.222
R3951 a_54966_3580.t0 a_54966_3580.t1 7.204
R3952 a_65700_25280.t0 a_65700_25280.t1 60
R3953 a_22972_23306.t0 a_22972_23306.n2 172.018
R3954 a_22972_23306.n2 a_22972_23306.t1 171.695
R3955 a_22972_23306.n2 a_22972_23306.n1 73.17
R3956 a_22972_23306.n1 a_22972_23306.t4 28.576
R3957 a_22972_23306.n0 a_22972_23306.t2 28.565
R3958 a_22972_23306.n0 a_22972_23306.t3 28.565
R3959 a_22972_23306.n1 a_22972_23306.n0 3.497
R3960 a_54468_7504.t0 a_54468_7504.t1 178.373
R3961 a_65689_26048.t0 a_65689_26048.t1 60
R3962 a_4314_11852.t0 a_4314_11852.t1 12.222
R3963 a_8748_11692.t0 a_8748_11692.t1 53.512
R3964 a_8748_9956.t0 a_8748_9956.t1 53.512
R3965 a_63985_26048.t1 a_63985_26048.t0 94.726
R3966 a_65523_26048.t0 a_65523_26048.t1 198.571
C19 vbiasot gnd 24.38fF $ **FLOATING
C20 vbiasob gnd 15.59fF $ **FLOATING
C21 z gnd 19.20fF $ **FLOATING
C22 vbiasbuffer gnd 16.94fF $ **FLOATING
C23 bb gnd 20.53fF $ **FLOATING
C24 aa gnd 22.72fF $ **FLOATING
C25 Fvco gnd 59.22fF $ **FLOATING
C26 vinit gnd 2.89fF $ **FLOATING
C27 Vso8b gnd 36.46fF $ **FLOATING
C28 Vso7b gnd 14.98fF $ **FLOATING
C29 Vso5b gnd 7.74fF $ **FLOATING
C30 Vso4b gnd 74.86fF $ **FLOATING
C31 Vso6b gnd 5.96fF $ **FLOATING
C32 vout gnd 8.80fF $ **FLOATING
C33 Fvco_By4_QPH_bar gnd 26.16fF $ **FLOATING
C34 Fvco_By4_QPH gnd 37.94fF $ **FLOATING
C35 RESET gnd 3.77fF $ **FLOATING
C36 CLK_IN gnd 46.25fF $ **FLOATING
C37 Vso3b gnd 45.20fF $ **FLOATING
C38 Vso2b gnd 33.81fF $ **FLOATING
C39 vctrl gnd 18.49fF $ **FLOATING
C40 zz gnd 5.84fF $ **FLOATING
C41 CLK_BY_4_IPH gnd 21.52fF
C42 CLK_BY_4_IPH_BAR gnd 69.13fF
C43 vdd gnd 5133.92fF
C44 a_54468_7504.t1 gnd 2.83fF
C45 a_22972_23306.n2 gnd 2.07fF $ **FLOATING
C46 a_47760_15642.n1 gnd 5.67fF $ **FLOATING
C47 a_47760_15642.n3 gnd 2.69fF $ **FLOATING
C48 a_42782_16060.n0 gnd 4.96fF $ **FLOATING
C49 a_42782_16060.n4 gnd 2.13fF $ **FLOATING
C50 a_43010_16058.n1 gnd 7.29fF $ **FLOATING
C51 a_43010_16058.n2 gnd 2.85fF $ **FLOATING
C52 Vso8b.n3 gnd 16.20fF $ **FLOATING
C53 a_4288_11726.n1 gnd 2.60fF $ **FLOATING
C54 a_4288_11726.n2 gnd 5.29fF $ **FLOATING
C55 aa.n3 gnd 8.25fF $ **FLOATING
C56 a_4226_11612.n1 gnd 4.10fF $ **FLOATING
C57 a_4226_11612.n2 gnd 5.11fF $ **FLOATING
C58 bb.n0 gnd 2.40fF $ **FLOATING
C59 bb.n11 gnd 8.77fF $ **FLOATING
C60 a_47968_16078.n0 gnd 4.32fF $ **FLOATING
C61 a_46856_19268.n0 gnd 7.50fF $ **FLOATING
C62 a_4288_12110.n1 gnd 4.71fF $ **FLOATING
C63 a_4288_12110.n2 gnd 3.47fF $ **FLOATING
C64 vbiasot.n1 gnd 6.96fF $ **FLOATING
C65 a_51138_21494.t0 gnd 2.55fF
C66 a_51138_21494.t1 gnd 3.48fF
C67 a_4226_11996.n1 gnd 4.19fF $ **FLOATING
C68 a_4226_11996.n2 gnd 6.64fF $ **FLOATING
C69 a_30384_802.n0 gnd 3.14fF $ **FLOATING
C70 a_38070_8852.n0 gnd 3.65fF $ **FLOATING
C71 a_50511_16072.n0 gnd 4.68fF $ **FLOATING
C72 a_50262_14152.n0 gnd 4.17fF $ **FLOATING
C73 a_51532_4150.n3 gnd 2.34fF $ **FLOATING
C74 a_51532_4150.n4 gnd 3.10fF $ **FLOATING
C75 a_4226_11804.n1 gnd 4.43fF $ **FLOATING
C76 a_4226_11804.n2 gnd 5.09fF $ **FLOATING
C77 Vso6b.n1 gnd 5.48fF $ **FLOATING
C78 Vso6b.n2 gnd 2.61fF $ **FLOATING
C79 z.n0 gnd 10.22fF $ **FLOATING
C80 a_51334_14126.n1 gnd 6.92fF $ **FLOATING
C81 Vso2b.n1 gnd 15.46fF $ **FLOATING
C82 a_28790_25040.n0 gnd 3.75fF $ **FLOATING
C83 a_32948_24994.n0 gnd 3.11fF $ **FLOATING
C84 a_4226_12188.n1 gnd 3.30fF $ **FLOATING
C85 a_4226_12188.n2 gnd 7.00fF $ **FLOATING
C86 a_23308_802.n0 gnd 3.31fF $ **FLOATING
C87 a_24410_25128.n0 gnd 3.81fF $ **FLOATING
C88 a_54448_7822.t0 gnd 3.00fF
C89 vout.n2 gnd 5.13fF $ **FLOATING
C90 a_4288_11918.n1 gnd 2.82fF $ **FLOATING
C91 a_4288_11918.n2 gnd 4.05fF $ **FLOATING
C92 Vso4b.n1 gnd 49.50fF $ **FLOATING
C93 a_14910_6932.n0 gnd 3.12fF $ **FLOATING
C94 a_42574_15624.n3 gnd 3.30fF $ **FLOATING
C95 a_42574_15624.n4 gnd 3.79fF $ **FLOATING
C96 a_42550_16062.n1 gnd 2.84fF $ **FLOATING
C97 a_42550_16062.n2 gnd 7.40fF $ **FLOATING
C98 Vso7b.n1 gnd 21.34fF $ **FLOATING
C99 Vso7b.n4 gnd 6.75fF $ **FLOATING
C100 CLK_BY_4_IPH_BAR.n2 gnd 2.98fF $ **FLOATING
C101 a_14832_12082.n0 gnd 3.86fF $ **FLOATING
C102 a_51138_19904.n0 gnd 2.56fF $ **FLOATING
C103 a_49932_4124.n1 gnd 2.10fF $ **FLOATING
C104 a_27762_11446.t21 gnd 11.67fF $ **FLOATING
C105 a_27762_11446.t11 gnd 33.06fF $ **FLOATING
C106 a_27762_11446.n0 gnd 3.93fF $ **FLOATING
C107 a_50583_13108.n0 gnd 8.05fF $ **FLOATING
C108 a_57726_5786.n0 gnd 2.08fF $ **FLOATING
C109 vbiasbuffer.n0 gnd 4.69fF $ **FLOATING
C110 vbiasob.n0 gnd 6.24fF $ **FLOATING
C111 a_56602_11692.n0 gnd 3.18fF $ **FLOATING
C112 Fvco.n0 gnd 4.49fF $ **FLOATING
C113 Fvco.n1 gnd 6.25fF $ **FLOATING
C114 Fvco.t34 gnd 2.57fF $ **FLOATING
C115 Fvco.n80 gnd 2.52fF $ **FLOATING
C116 Fvco.n81 gnd 38.82fF $ **FLOATING
C117 a_4288_11534.n1 gnd 2.34fF $ **FLOATING
C118 a_4288_11534.n2 gnd 4.20fF $ **FLOATING
C119 CLK_IN.n0 gnd 2.40fF $ **FLOATING
C120 CLK_IN.n1 gnd 46.02fF $ **FLOATING
C121 CLK_IN.n4 gnd 12.12fF $ **FLOATING
C122 a_51276_14152.n1 gnd 3.79fF $ **FLOATING
C123 a_51636_13108.n3 gnd 2.84fF $ **FLOATING
C124 a_23436_16644.t12 gnd 32.42fF $ **FLOATING
C125 a_23436_16644.n0 gnd 3.27fF $ **FLOATING
C126 a_56334_20860.n0 gnd 2.57fF $ **FLOATING
C127 a_52052_20860.t0 gnd 3.50fF
C128 Vso5b.n1 gnd 8.15fF $ **FLOATING
C129 Vso5b.n2 gnd 3.73fF $ **FLOATING
C130 Vso3b.n1 gnd 11.41fF $ **FLOATING
C131 a_14266_8900.t47 gnd 27.25fF $ **FLOATING
C132 a_14266_8900.t16 gnd 23.08fF $ **FLOATING
C133 a_17685_3840.t22 gnd 2.79fF $ **FLOATING
C134 a_17685_3840.t63 gnd 2.79fF $ **FLOATING
C135 a_17685_3840.t58 gnd 2.79fF $ **FLOATING
C136 a_17685_3840.t60 gnd 2.79fF $ **FLOATING
C137 a_17685_3840.t53 gnd 2.79fF $ **FLOATING
C138 a_17685_3840.t48 gnd 2.79fF $ **FLOATING
C139 a_17685_3840.t20 gnd 2.79fF $ **FLOATING
C140 a_17685_3840.t64 gnd 2.79fF $ **FLOATING
C141 a_17685_3840.t56 gnd 2.79fF $ **FLOATING
C142 a_17685_3840.t51 gnd 2.79fF $ **FLOATING
C143 a_17685_3840.t43 gnd 6.44fF $ **FLOATING
C144 a_17685_3840.n1 gnd 11.37fF $ **FLOATING
C145 a_17685_3840.n2 gnd 7.40fF $ **FLOATING
C146 a_17685_3840.n3 gnd 7.40fF $ **FLOATING
C147 a_17685_3840.n4 gnd 7.40fF $ **FLOATING
C148 a_17685_3840.n5 gnd 7.40fF $ **FLOATING
C149 a_17685_3840.n6 gnd 7.40fF $ **FLOATING
C150 a_17685_3840.n7 gnd 7.40fF $ **FLOATING
C151 a_17685_3840.n8 gnd 7.40fF $ **FLOATING
C152 a_17685_3840.n9 gnd 7.40fF $ **FLOATING
C153 a_17685_3840.n10 gnd 6.25fF $ **FLOATING
C154 a_17685_3840.t54 gnd 3.74fF $ **FLOATING
C155 a_17685_3840.n11 gnd 7.66fF $ **FLOATING
C156 a_17685_3840.t46 gnd 2.79fF $ **FLOATING
C157 a_17685_3840.t38 gnd 2.79fF $ **FLOATING
C158 a_17685_3840.t31 gnd 2.79fF $ **FLOATING
C159 a_17685_3840.t33 gnd 2.79fF $ **FLOATING
C160 a_17685_3840.t24 gnd 2.79fF $ **FLOATING
C161 a_17685_3840.t18 gnd 2.79fF $ **FLOATING
C162 a_17685_3840.t61 gnd 2.79fF $ **FLOATING
C163 a_17685_3840.t55 gnd 2.79fF $ **FLOATING
C164 a_17685_3840.t49 gnd 2.79fF $ **FLOATING
C165 a_17685_3840.t42 gnd 2.79fF $ **FLOATING
C166 a_17685_3840.t35 gnd 6.44fF $ **FLOATING
C167 a_17685_3840.n12 gnd 11.34fF $ **FLOATING
C168 a_17685_3840.n13 gnd 7.39fF $ **FLOATING
C169 a_17685_3840.n14 gnd 7.39fF $ **FLOATING
C170 a_17685_3840.n15 gnd 7.39fF $ **FLOATING
C171 a_17685_3840.n16 gnd 7.39fF $ **FLOATING
C172 a_17685_3840.n17 gnd 7.39fF $ **FLOATING
C173 a_17685_3840.n18 gnd 7.39fF $ **FLOATING
C174 a_17685_3840.n19 gnd 7.39fF $ **FLOATING
C175 a_17685_3840.n20 gnd 7.39fF $ **FLOATING
C176 a_17685_3840.n21 gnd 6.25fF $ **FLOATING
C177 a_17685_3840.t27 gnd 3.74fF $ **FLOATING
C178 a_17685_3840.n22 gnd 5.61fF $ **FLOATING
C179 a_17685_3840.n23 gnd 6.37fF $ **FLOATING
C180 a_17685_3840.n24 gnd 3.21fF $ **FLOATING
C181 a_17685_3840.n29 gnd 2.54fF $ **FLOATING
C182 a_17685_3840.t47 gnd 2.79fF $ **FLOATING
C183 a_17685_3840.t41 gnd 2.79fF $ **FLOATING
C184 a_17685_3840.t44 gnd 2.79fF $ **FLOATING
C185 a_17685_3840.t36 gnd 2.79fF $ **FLOATING
C186 a_17685_3840.t29 gnd 2.79fF $ **FLOATING
C187 a_17685_3840.t28 gnd 2.79fF $ **FLOATING
C188 a_17685_3840.t21 gnd 2.79fF $ **FLOATING
C189 a_17685_3840.t62 gnd 2.79fF $ **FLOATING
C190 a_17685_3840.t57 gnd 2.79fF $ **FLOATING
C191 a_17685_3840.t50 gnd 6.44fF $ **FLOATING
C192 a_17685_3840.n34 gnd 11.33fF $ **FLOATING
C193 a_17685_3840.n35 gnd 7.38fF $ **FLOATING
C194 a_17685_3840.n36 gnd 7.38fF $ **FLOATING
C195 a_17685_3840.n37 gnd 7.38fF $ **FLOATING
C196 a_17685_3840.n38 gnd 7.38fF $ **FLOATING
C197 a_17685_3840.n39 gnd 7.38fF $ **FLOATING
C198 a_17685_3840.n40 gnd 7.38fF $ **FLOATING
C199 a_17685_3840.n41 gnd 7.38fF $ **FLOATING
C200 a_17685_3840.n42 gnd 7.38fF $ **FLOATING
C201 a_17685_3840.t52 gnd 2.79fF $ **FLOATING
C202 a_17685_3840.n43 gnd 6.22fF $ **FLOATING
C203 a_17685_3840.t39 gnd 3.75fF $ **FLOATING
C204 a_17685_3840.n44 gnd 7.71fF $ **FLOATING
C205 a_17685_3840.t45 gnd 2.79fF $ **FLOATING
C206 a_17685_3840.t37 gnd 2.79fF $ **FLOATING
C207 a_17685_3840.t30 gnd 2.79fF $ **FLOATING
C208 a_17685_3840.t32 gnd 2.79fF $ **FLOATING
C209 a_17685_3840.t23 gnd 2.79fF $ **FLOATING
C210 a_17685_3840.t17 gnd 2.79fF $ **FLOATING
C211 a_17685_3840.t40 gnd 2.79fF $ **FLOATING
C212 a_17685_3840.t34 gnd 2.79fF $ **FLOATING
C213 a_17685_3840.t25 gnd 2.79fF $ **FLOATING
C214 a_17685_3840.t19 gnd 2.79fF $ **FLOATING
C215 a_17685_3840.t59 gnd 6.45fF $ **FLOATING
C216 a_17685_3840.n45 gnd 11.38fF $ **FLOATING
C217 a_17685_3840.n46 gnd 7.41fF $ **FLOATING
C218 a_17685_3840.n47 gnd 7.41fF $ **FLOATING
C219 a_17685_3840.n48 gnd 7.41fF $ **FLOATING
C220 a_17685_3840.n49 gnd 7.41fF $ **FLOATING
C221 a_17685_3840.n50 gnd 7.41fF $ **FLOATING
C222 a_17685_3840.n51 gnd 7.41fF $ **FLOATING
C223 a_17685_3840.n52 gnd 7.41fF $ **FLOATING
C224 a_17685_3840.n53 gnd 7.41fF $ **FLOATING
C225 a_17685_3840.n54 gnd 6.26fF $ **FLOATING
C226 a_17685_3840.t26 gnd 3.74fF $ **FLOATING
C227 a_17685_3840.n55 gnd 5.44fF $ **FLOATING
C228 a_17685_3840.n56 gnd 6.26fF $ **FLOATING
C229 a_17685_3840.n57 gnd 3.40fF $ **FLOATING
C230 a_17685_3840.n60 gnd 2.24fF $ **FLOATING
C231 a_25099_11445.t15 gnd 26.39fF $ **FLOATING
C232 a_25099_11445.t52 gnd 18.22fF $ **FLOATING
C233 vctrl.n2 gnd 5.05fF $ **FLOATING
C234 CLK_BY_4_IPH.n3 gnd 29.42fF $ **FLOATING
C235 a_26036_4988.t20 gnd 21.24fF $ **FLOATING
C236 a_26036_4988.t16 gnd 15.27fF $ **FLOATING
C237 a_14188_14050.t31 gnd 36.88fF $ **FLOATING
C238 a_14188_14050.t12 gnd 24.22fF $ **FLOATING
C239 a_49874_4150.t0 gnd 11.61fF
C240 a_49874_4150.t1 gnd 9.04fF
C241 a_50320_14126.n6 gnd 8.78fF $ **FLOATING
C242 a_50320_14126.n7 gnd 2.15fF $ **FLOATING
C243 a_55602_11692.n0 gnd 2.80fF $ **FLOATING
C244 Fvco_By4_QPH.n0 gnd 11.76fF $ **FLOATING
C245 Fvco_By4_QPH.n2 gnd 2.48fF $ **FLOATING
C246 Fvco_By4_QPH.n3 gnd 2.45fF $ **FLOATING
C247 Fvco_By4_QPH.n4 gnd 5.17fF $ **FLOATING
C248 Fvco_By4_QPH.n6 gnd 5.63fF $ **FLOATING
C249 a_4226_11420.n1 gnd 3.51fF $ **FLOATING
C250 a_4226_11420.n2 gnd 5.45fF $ **FLOATING
C251 Vso1b.n0 gnd 20.26fF $ **FLOATING
C252 Vso1b.n3 gnd 12.35fF $ **FLOATING
C253 a_1026_45630.t73 gnd 6.88fF $ **FLOATING
C254 a_1026_45630.n2 gnd 8.73fF $ **FLOATING
C255 a_1026_45630.t7 gnd 2.37fF $ **FLOATING
C256 a_1026_45630.n3 gnd 6.45fF $ **FLOATING
C257 a_1026_45630.t44 gnd 2.37fF $ **FLOATING
C258 a_1026_45630.n4 gnd 6.33fF $ **FLOATING
C259 a_1026_45630.t202 gnd 2.37fF $ **FLOATING
C260 a_1026_45630.n5 gnd 6.33fF $ **FLOATING
C261 a_1026_45630.t133 gnd 2.37fF $ **FLOATING
C262 a_1026_45630.n6 gnd 6.33fF $ **FLOATING
C263 a_1026_45630.t180 gnd 2.37fF $ **FLOATING
C264 a_1026_45630.n7 gnd 6.33fF $ **FLOATING
C265 a_1026_45630.t129 gnd 2.37fF $ **FLOATING
C266 a_1026_45630.n8 gnd 6.33fF $ **FLOATING
C267 a_1026_45630.t59 gnd 2.37fF $ **FLOATING
C268 a_1026_45630.n9 gnd 6.33fF $ **FLOATING
C269 a_1026_45630.t18 gnd 2.37fF $ **FLOATING
C270 a_1026_45630.n10 gnd 3.52fF $ **FLOATING
C271 a_1026_45630.t147 gnd 2.37fF $ **FLOATING
C272 a_1026_45630.t172 gnd 6.85fF $ **FLOATING
C273 a_1026_45630.n11 gnd 8.72fF $ **FLOATING
C274 a_1026_45630.t105 gnd 2.37fF $ **FLOATING
C275 a_1026_45630.n12 gnd 6.45fF $ **FLOATING
C276 a_1026_45630.t190 gnd 2.37fF $ **FLOATING
C277 a_1026_45630.n13 gnd 6.33fF $ **FLOATING
C278 a_1026_45630.t143 gnd 2.37fF $ **FLOATING
C279 a_1026_45630.n14 gnd 6.33fF $ **FLOATING
C280 a_1026_45630.t76 gnd 2.37fF $ **FLOATING
C281 a_1026_45630.n15 gnd 6.33fF $ **FLOATING
C282 a_1026_45630.t123 gnd 2.37fF $ **FLOATING
C283 a_1026_45630.n16 gnd 6.33fF $ **FLOATING
C284 a_1026_45630.t72 gnd 2.37fF $ **FLOATING
C285 a_1026_45630.n17 gnd 6.33fF $ **FLOATING
C286 a_1026_45630.t6 gnd 2.37fF $ **FLOATING
C287 a_1026_45630.n18 gnd 6.33fF $ **FLOATING
C288 a_1026_45630.t159 gnd 2.37fF $ **FLOATING
C289 a_1026_45630.n19 gnd 3.36fF $ **FLOATING
C290 a_1026_45630.t96 gnd 2.37fF $ **FLOATING
C291 a_1026_45630.n20 gnd 6.33fF $ **FLOATING
C292 a_1026_45630.t138 gnd 2.37fF $ **FLOATING
C293 a_1026_45630.n21 gnd 6.33fF $ **FLOATING
C294 a_1026_45630.t5 gnd 2.37fF $ **FLOATING
C295 a_1026_45630.n22 gnd 6.33fF $ **FLOATING
C296 a_1026_45630.t48 gnd 2.37fF $ **FLOATING
C297 a_1026_45630.n23 gnd 6.33fF $ **FLOATING
C298 a_1026_45630.t117 gnd 2.37fF $ **FLOATING
C299 a_1026_45630.n24 gnd 6.33fF $ **FLOATING
C300 a_1026_45630.t170 gnd 2.37fF $ **FLOATING
C301 a_1026_45630.n25 gnd 6.33fF $ **FLOATING
C302 a_1026_45630.t121 gnd 2.37fF $ **FLOATING
C303 a_1026_45630.n26 gnd 6.33fF $ **FLOATING
C304 a_1026_45630.t188 gnd 2.37fF $ **FLOATING
C305 a_1026_45630.n27 gnd 6.45fF $ **FLOATING
C306 a_1026_45630.t33 gnd 2.37fF $ **FLOATING
C307 a_1026_45630.n28 gnd 8.69fF $ **FLOATING
C308 a_1026_45630.t148 gnd 2.37fF $ **FLOATING
C309 a_1026_45630.t17 gnd 6.78fF $ **FLOATING
C310 a_1026_45630.n29 gnd 3.03fF $ **FLOATING
C311 a_1026_45630.t131 gnd 6.88fF $ **FLOATING
C312 a_1026_45630.n30 gnd 8.73fF $ **FLOATING
C313 a_1026_45630.t60 gnd 2.37fF $ **FLOATING
C314 a_1026_45630.n31 gnd 6.45fF $ **FLOATING
C315 a_1026_45630.t150 gnd 2.37fF $ **FLOATING
C316 a_1026_45630.n32 gnd 6.33fF $ **FLOATING
C317 a_1026_45630.t107 gnd 2.37fF $ **FLOATING
C318 a_1026_45630.n33 gnd 6.33fF $ **FLOATING
C319 a_1026_45630.t34 gnd 2.37fF $ **FLOATING
C320 a_1026_45630.n34 gnd 6.33fF $ **FLOATING
C321 a_1026_45630.t85 gnd 2.37fF $ **FLOATING
C322 a_1026_45630.n35 gnd 6.33fF $ **FLOATING
C323 a_1026_45630.t30 gnd 2.37fF $ **FLOATING
C324 a_1026_45630.n36 gnd 6.33fF $ **FLOATING
C325 a_1026_45630.t163 gnd 2.37fF $ **FLOATING
C326 a_1026_45630.n37 gnd 6.33fF $ **FLOATING
C327 a_1026_45630.t118 gnd 2.37fF $ **FLOATING
C328 a_1026_45630.n38 gnd 3.52fF $ **FLOATING
C329 a_1026_45630.t49 gnd 2.37fF $ **FLOATING
C330 a_1026_45630.n39 gnd 2.93fF $ **FLOATING
C331 a_1026_45630.t95 gnd 6.78fF $ **FLOATING
C332 a_1026_45630.n40 gnd 8.69fF $ **FLOATING
C333 a_1026_45630.t24 gnd 2.37fF $ **FLOATING
C334 a_1026_45630.n41 gnd 6.45fF $ **FLOATING
C335 a_1026_45630.t112 gnd 2.37fF $ **FLOATING
C336 a_1026_45630.n42 gnd 6.33fF $ **FLOATING
C337 a_1026_45630.t64 gnd 2.37fF $ **FLOATING
C338 a_1026_45630.n43 gnd 6.33fF $ **FLOATING
C339 a_1026_45630.t195 gnd 2.37fF $ **FLOATING
C340 a_1026_45630.n44 gnd 6.33fF $ **FLOATING
C341 a_1026_45630.t43 gnd 2.37fF $ **FLOATING
C342 a_1026_45630.n45 gnd 6.33fF $ **FLOATING
C343 a_1026_45630.t191 gnd 2.37fF $ **FLOATING
C344 a_1026_45630.n46 gnd 6.33fF $ **FLOATING
C345 a_1026_45630.t124 gnd 2.37fF $ **FLOATING
C346 a_1026_45630.n47 gnd 6.33fF $ **FLOATING
C347 a_1026_45630.t77 gnd 2.37fF $ **FLOATING
C348 a_1026_45630.n48 gnd 3.52fF $ **FLOATING
C349 a_1026_45630.t12 gnd 2.37fF $ **FLOATING
C350 a_1026_45630.n49 gnd 2.94fF $ **FLOATING
C351 a_1026_45630.t45 gnd 6.88fF $ **FLOATING
C352 a_1026_45630.n50 gnd 8.73fF $ **FLOATING
C353 a_1026_45630.t182 gnd 2.37fF $ **FLOATING
C354 a_1026_45630.n51 gnd 6.45fF $ **FLOATING
C355 a_1026_45630.t70 gnd 2.37fF $ **FLOATING
C356 a_1026_45630.n52 gnd 6.33fF $ **FLOATING
C357 a_1026_45630.t26 gnd 2.37fF $ **FLOATING
C358 a_1026_45630.n53 gnd 6.33fF $ **FLOATING
C359 a_1026_45630.t157 gnd 2.37fF $ **FLOATING
C360 a_1026_45630.n54 gnd 6.33fF $ **FLOATING
C361 a_1026_45630.t4 gnd 2.37fF $ **FLOATING
C362 a_1026_45630.n55 gnd 6.33fF $ **FLOATING
C363 a_1026_45630.t153 gnd 2.37fF $ **FLOATING
C364 a_1026_45630.n56 gnd 6.33fF $ **FLOATING
C365 a_1026_45630.t87 gnd 2.37fF $ **FLOATING
C366 a_1026_45630.n57 gnd 6.33fF $ **FLOATING
C367 a_1026_45630.t37 gnd 2.37fF $ **FLOATING
C368 a_1026_45630.n58 gnd 3.52fF $ **FLOATING
C369 a_1026_45630.t173 gnd 2.37fF $ **FLOATING
C370 a_1026_45630.n59 gnd 2.93fF $ **FLOATING
C371 a_1026_45630.t15 gnd 6.85fF $ **FLOATING
C372 a_1026_45630.n60 gnd 8.72fF $ **FLOATING
C373 a_1026_45630.t144 gnd 2.37fF $ **FLOATING
C374 a_1026_45630.n61 gnd 6.45fF $ **FLOATING
C375 a_1026_45630.t184 gnd 2.37fF $ **FLOATING
C376 a_1026_45630.n62 gnd 6.33fF $ **FLOATING
C377 a_1026_45630.t139 gnd 2.37fF $ **FLOATING
C378 a_1026_45630.n63 gnd 6.33fF $ **FLOATING
C379 a_1026_45630.t71 gnd 2.37fF $ **FLOATING
C380 a_1026_45630.n64 gnd 6.33fF $ **FLOATING
C381 a_1026_45630.t116 gnd 2.37fF $ **FLOATING
C382 a_1026_45630.n65 gnd 6.33fF $ **FLOATING
C383 a_1026_45630.t67 gnd 2.37fF $ **FLOATING
C384 a_1026_45630.n66 gnd 6.33fF $ **FLOATING
C385 a_1026_45630.t201 gnd 2.37fF $ **FLOATING
C386 a_1026_45630.n67 gnd 6.33fF $ **FLOATING
C387 a_1026_45630.t155 gnd 2.37fF $ **FLOATING
C388 a_1026_45630.n68 gnd 3.52fF $ **FLOATING
C389 a_1026_45630.t89 gnd 2.37fF $ **FLOATING
C390 a_1026_45630.n69 gnd 2.94fF $ **FLOATING
C391 a_1026_45630.t177 gnd 6.88fF $ **FLOATING
C392 a_1026_45630.n70 gnd 8.73fF $ **FLOATING
C393 a_1026_45630.t109 gnd 2.37fF $ **FLOATING
C394 a_1026_45630.n71 gnd 6.45fF $ **FLOATING
C395 a_1026_45630.t193 gnd 2.37fF $ **FLOATING
C396 a_1026_45630.n72 gnd 6.33fF $ **FLOATING
C397 a_1026_45630.t149 gnd 2.37fF $ **FLOATING
C398 a_1026_45630.n73 gnd 6.33fF $ **FLOATING
C399 a_1026_45630.t79 gnd 2.37fF $ **FLOATING
C400 a_1026_45630.n74 gnd 6.33fF $ **FLOATING
C401 a_1026_45630.t128 gnd 2.37fF $ **FLOATING
C402 a_1026_45630.n75 gnd 6.33fF $ **FLOATING
C403 a_1026_45630.t75 gnd 2.37fF $ **FLOATING
C404 a_1026_45630.n76 gnd 6.33fF $ **FLOATING
C405 a_1026_45630.t8 gnd 2.37fF $ **FLOATING
C406 a_1026_45630.n77 gnd 6.33fF $ **FLOATING
C407 a_1026_45630.t161 gnd 2.37fF $ **FLOATING
C408 a_1026_45630.n78 gnd 3.52fF $ **FLOATING
C409 a_1026_45630.t98 gnd 2.37fF $ **FLOATING
C410 a_1026_45630.n79 gnd 2.93fF $ **FLOATING
C411 a_1026_45630.t127 gnd 6.82fF $ **FLOATING
C412 a_1026_45630.n80 gnd 8.70fF $ **FLOATING
C413 a_1026_45630.t56 gnd 2.37fF $ **FLOATING
C414 a_1026_45630.n81 gnd 6.45fF $ **FLOATING
C415 a_1026_45630.t146 gnd 2.37fF $ **FLOATING
C416 a_1026_45630.n82 gnd 6.33fF $ **FLOATING
C417 a_1026_45630.t102 gnd 2.37fF $ **FLOATING
C418 a_1026_45630.n83 gnd 6.33fF $ **FLOATING
C419 a_1026_45630.t32 gnd 2.37fF $ **FLOATING
C420 a_1026_45630.n84 gnd 6.33fF $ **FLOATING
C421 a_1026_45630.t81 gnd 2.37fF $ **FLOATING
C422 a_1026_45630.n85 gnd 6.33fF $ **FLOATING
C423 a_1026_45630.t28 gnd 2.37fF $ **FLOATING
C424 a_1026_45630.n86 gnd 6.33fF $ **FLOATING
C425 a_1026_45630.t160 gnd 2.37fF $ **FLOATING
C426 a_1026_45630.n87 gnd 6.33fF $ **FLOATING
C427 a_1026_45630.t115 gnd 2.37fF $ **FLOATING
C428 a_1026_45630.n88 gnd 3.52fF $ **FLOATING
C429 a_1026_45630.t46 gnd 2.37fF $ **FLOATING
C430 a_1026_45630.n89 gnd 2.93fF $ **FLOATING
C431 a_1026_45630.t91 gnd 6.85fF $ **FLOATING
C432 a_1026_45630.n90 gnd 8.72fF $ **FLOATING
C433 a_1026_45630.t21 gnd 2.37fF $ **FLOATING
C434 a_1026_45630.n91 gnd 6.45fF $ **FLOATING
C435 a_1026_45630.t111 gnd 2.37fF $ **FLOATING
C436 a_1026_45630.n92 gnd 6.33fF $ **FLOATING
C437 a_1026_45630.t58 gnd 2.37fF $ **FLOATING
C438 a_1026_45630.n93 gnd 6.33fF $ **FLOATING
C439 a_1026_45630.t192 gnd 2.37fF $ **FLOATING
C440 a_1026_45630.n94 gnd 6.33fF $ **FLOATING
C441 a_1026_45630.t41 gnd 2.37fF $ **FLOATING
C442 a_1026_45630.n95 gnd 6.33fF $ **FLOATING
C443 a_1026_45630.t189 gnd 2.37fF $ **FLOATING
C444 a_1026_45630.n96 gnd 6.33fF $ **FLOATING
C445 a_1026_45630.t122 gnd 2.37fF $ **FLOATING
C446 a_1026_45630.n97 gnd 6.33fF $ **FLOATING
C447 a_1026_45630.t74 gnd 2.37fF $ **FLOATING
C448 a_1026_45630.n98 gnd 3.52fF $ **FLOATING
C449 a_1026_45630.t9 gnd 2.37fF $ **FLOATING
C450 a_1026_45630.n99 gnd 2.94fF $ **FLOATING
C451 a_1026_45630.t179 gnd 6.82fF $ **FLOATING
C452 a_1026_45630.n100 gnd 8.70fF $ **FLOATING
C453 a_1026_45630.t113 gnd 2.37fF $ **FLOATING
C454 a_1026_45630.n101 gnd 6.45fF $ **FLOATING
C455 a_1026_45630.t200 gnd 2.37fF $ **FLOATING
C456 a_1026_45630.n102 gnd 6.33fF $ **FLOATING
C457 a_1026_45630.t154 gnd 2.37fF $ **FLOATING
C458 a_1026_45630.n103 gnd 6.33fF $ **FLOATING
C459 a_1026_45630.t90 gnd 2.37fF $ **FLOATING
C460 a_1026_45630.n104 gnd 6.33fF $ **FLOATING
C461 a_1026_45630.t134 gnd 2.37fF $ **FLOATING
C462 a_1026_45630.n105 gnd 6.33fF $ **FLOATING
C463 a_1026_45630.t82 gnd 2.37fF $ **FLOATING
C464 a_1026_45630.n106 gnd 6.33fF $ **FLOATING
C465 a_1026_45630.t16 gnd 2.37fF $ **FLOATING
C466 a_1026_45630.n107 gnd 6.33fF $ **FLOATING
C467 a_1026_45630.t167 gnd 2.37fF $ **FLOATING
C468 a_1026_45630.n108 gnd 3.52fF $ **FLOATING
C469 a_1026_45630.t101 gnd 2.37fF $ **FLOATING
C470 a_1026_45630.n109 gnd 2.93fF $ **FLOATING
C471 a_1026_45630.t11 gnd 6.85fF $ **FLOATING
C472 a_1026_45630.n110 gnd 8.72fF $ **FLOATING
C473 a_1026_45630.t141 gnd 2.37fF $ **FLOATING
C474 a_1026_45630.n111 gnd 6.45fF $ **FLOATING
C475 a_1026_45630.t181 gnd 2.37fF $ **FLOATING
C476 a_1026_45630.n112 gnd 6.33fF $ **FLOATING
C477 a_1026_45630.t135 gnd 2.37fF $ **FLOATING
C478 a_1026_45630.n113 gnd 6.33fF $ **FLOATING
C479 a_1026_45630.t68 gnd 2.37fF $ **FLOATING
C480 a_1026_45630.n114 gnd 6.33fF $ **FLOATING
C481 a_1026_45630.t114 gnd 2.37fF $ **FLOATING
C482 a_1026_45630.n115 gnd 6.33fF $ **FLOATING
C483 a_1026_45630.t63 gnd 2.37fF $ **FLOATING
C484 a_1026_45630.n116 gnd 6.33fF $ **FLOATING
C485 a_1026_45630.t196 gnd 2.37fF $ **FLOATING
C486 a_1026_45630.n117 gnd 6.33fF $ **FLOATING
C487 a_1026_45630.t151 gnd 2.37fF $ **FLOATING
C488 a_1026_45630.n118 gnd 3.52fF $ **FLOATING
C489 a_1026_45630.t83 gnd 2.37fF $ **FLOATING
C490 a_1026_45630.n119 gnd 3.09fF $ **FLOATING
C491 a_1026_45630.n120 gnd 2.94fF $ **FLOATING
C492 a_1026_45630.t61 gnd 6.88fF $ **FLOATING
C493 a_1026_45630.n121 gnd 8.73fF $ **FLOATING
C494 a_1026_45630.t194 gnd 2.37fF $ **FLOATING
C495 a_1026_45630.n122 gnd 6.45fF $ **FLOATING
C496 a_1026_45630.t84 gnd 2.37fF $ **FLOATING
C497 a_1026_45630.n123 gnd 6.33fF $ **FLOATING
C498 a_1026_45630.t35 gnd 2.37fF $ **FLOATING
C499 a_1026_45630.n124 gnd 6.33fF $ **FLOATING
C500 a_1026_45630.t171 gnd 2.37fF $ **FLOATING
C501 a_1026_45630.n125 gnd 6.33fF $ **FLOATING
C502 a_1026_45630.t19 gnd 2.37fF $ **FLOATING
C503 a_1026_45630.n126 gnd 6.33fF $ **FLOATING
C504 a_1026_45630.t164 gnd 2.37fF $ **FLOATING
C505 a_1026_45630.n127 gnd 6.33fF $ **FLOATING
C506 a_1026_45630.t99 gnd 2.37fF $ **FLOATING
C507 a_1026_45630.n128 gnd 6.33fF $ **FLOATING
C508 a_1026_45630.t50 gnd 2.37fF $ **FLOATING
C509 a_1026_45630.n129 gnd 3.52fF $ **FLOATING
C510 a_1026_45630.t185 gnd 2.37fF $ **FLOATING
C511 a_1026_45630.n130 gnd 2.93fF $ **FLOATING
C512 a_1026_45630.t132 gnd 6.88fF $ **FLOATING
C513 a_1026_45630.n131 gnd 8.73fF $ **FLOATING
C514 a_1026_45630.t62 gnd 2.37fF $ **FLOATING
C515 a_1026_45630.n132 gnd 6.45fF $ **FLOATING
C516 a_1026_45630.t152 gnd 2.37fF $ **FLOATING
C517 a_1026_45630.n133 gnd 6.33fF $ **FLOATING
C518 a_1026_45630.t108 gnd 2.37fF $ **FLOATING
C519 a_1026_45630.n134 gnd 6.33fF $ **FLOATING
C520 a_1026_45630.t36 gnd 2.37fF $ **FLOATING
C521 a_1026_45630.n135 gnd 6.33fF $ **FLOATING
C522 a_1026_45630.t86 gnd 2.37fF $ **FLOATING
C523 a_1026_45630.n136 gnd 6.33fF $ **FLOATING
C524 a_1026_45630.t31 gnd 2.37fF $ **FLOATING
C525 a_1026_45630.n137 gnd 6.33fF $ **FLOATING
C526 a_1026_45630.t165 gnd 2.37fF $ **FLOATING
C527 a_1026_45630.n138 gnd 6.33fF $ **FLOATING
C528 a_1026_45630.t119 gnd 2.37fF $ **FLOATING
C529 a_1026_45630.n139 gnd 3.52fF $ **FLOATING
C530 a_1026_45630.t51 gnd 2.37fF $ **FLOATING
C531 a_1026_45630.n140 gnd 2.93fF $ **FLOATING
C532 a_1026_45630.t25 gnd 6.88fF $ **FLOATING
C533 a_1026_45630.n141 gnd 8.73fF $ **FLOATING
C534 a_1026_45630.t156 gnd 2.37fF $ **FLOATING
C535 a_1026_45630.n142 gnd 6.45fF $ **FLOATING
C536 a_1026_45630.t42 gnd 2.37fF $ **FLOATING
C537 a_1026_45630.n143 gnd 6.33fF $ **FLOATING
C538 a_1026_45630.t197 gnd 2.37fF $ **FLOATING
C539 a_1026_45630.n144 gnd 6.33fF $ **FLOATING
C540 a_1026_45630.t130 gnd 2.37fF $ **FLOATING
C541 a_1026_45630.n145 gnd 6.33fF $ **FLOATING
C542 a_1026_45630.t178 gnd 2.37fF $ **FLOATING
C543 a_1026_45630.n146 gnd 6.33fF $ **FLOATING
C544 a_1026_45630.t125 gnd 2.37fF $ **FLOATING
C545 a_1026_45630.n147 gnd 6.33fF $ **FLOATING
C546 a_1026_45630.t55 gnd 2.37fF $ **FLOATING
C547 a_1026_45630.n148 gnd 6.33fF $ **FLOATING
C548 a_1026_45630.t13 gnd 2.37fF $ **FLOATING
C549 a_1026_45630.n149 gnd 3.52fF $ **FLOATING
C550 a_1026_45630.t142 gnd 2.37fF $ **FLOATING
C551 a_1026_45630.n150 gnd 2.94fF $ **FLOATING
C552 a_1026_45630.t29 gnd 6.88fF $ **FLOATING
C553 a_1026_45630.n151 gnd 8.73fF $ **FLOATING
C554 a_1026_45630.t162 gnd 2.37fF $ **FLOATING
C555 a_1026_45630.n152 gnd 6.45fF $ **FLOATING
C556 a_1026_45630.t203 gnd 2.37fF $ **FLOATING
C557 a_1026_45630.n153 gnd 6.33fF $ **FLOATING
C558 a_1026_45630.t158 gnd 2.37fF $ **FLOATING
C559 a_1026_45630.n154 gnd 6.33fF $ **FLOATING
C560 a_1026_45630.t94 gnd 2.37fF $ **FLOATING
C561 a_1026_45630.n155 gnd 6.33fF $ **FLOATING
C562 a_1026_45630.t136 gnd 2.37fF $ **FLOATING
C563 a_1026_45630.n156 gnd 6.33fF $ **FLOATING
C564 a_1026_45630.t88 gnd 2.37fF $ **FLOATING
C565 a_1026_45630.n157 gnd 6.33fF $ **FLOATING
C566 a_1026_45630.t20 gnd 2.37fF $ **FLOATING
C567 a_1026_45630.n158 gnd 6.33fF $ **FLOATING
C568 a_1026_45630.t174 gnd 2.37fF $ **FLOATING
C569 a_1026_45630.n159 gnd 3.52fF $ **FLOATING
C570 a_1026_45630.t106 gnd 2.37fF $ **FLOATING
C571 a_1026_45630.n160 gnd 2.94fF $ **FLOATING
C572 a_1026_45630.t145 gnd 6.85fF $ **FLOATING
C573 a_1026_45630.n161 gnd 8.72fF $ **FLOATING
C574 a_1026_45630.t78 gnd 2.37fF $ **FLOATING
C575 a_1026_45630.n162 gnd 6.45fF $ **FLOATING
C576 a_1026_45630.t166 gnd 2.37fF $ **FLOATING
C577 a_1026_45630.n163 gnd 6.33fF $ **FLOATING
C578 a_1026_45630.t120 gnd 2.37fF $ **FLOATING
C579 a_1026_45630.n164 gnd 6.33fF $ **FLOATING
C580 a_1026_45630.t52 gnd 2.37fF $ **FLOATING
C581 a_1026_45630.n165 gnd 6.33fF $ **FLOATING
C582 a_1026_45630.t100 gnd 2.37fF $ **FLOATING
C583 a_1026_45630.n166 gnd 6.33fF $ **FLOATING
C584 a_1026_45630.t47 gnd 2.37fF $ **FLOATING
C585 a_1026_45630.n167 gnd 6.33fF $ **FLOATING
C586 a_1026_45630.t183 gnd 2.37fF $ **FLOATING
C587 a_1026_45630.n168 gnd 6.33fF $ **FLOATING
C588 a_1026_45630.t137 gnd 2.37fF $ **FLOATING
C589 a_1026_45630.n169 gnd 3.52fF $ **FLOATING
C590 a_1026_45630.t69 gnd 2.37fF $ **FLOATING
C591 a_1026_45630.n170 gnd 2.93fF $ **FLOATING
C592 a_1026_45630.t110 gnd 6.91fF $ **FLOATING
C593 a_1026_45630.n171 gnd 8.75fF $ **FLOATING
C594 a_1026_45630.t38 gnd 2.37fF $ **FLOATING
C595 a_1026_45630.n172 gnd 6.45fF $ **FLOATING
C596 a_1026_45630.t126 gnd 2.37fF $ **FLOATING
C597 a_1026_45630.n173 gnd 6.33fF $ **FLOATING
C598 a_1026_45630.t80 gnd 2.37fF $ **FLOATING
C599 a_1026_45630.n174 gnd 6.33fF $ **FLOATING
C600 a_1026_45630.t14 gnd 2.37fF $ **FLOATING
C601 a_1026_45630.n175 gnd 6.33fF $ **FLOATING
C602 a_1026_45630.t57 gnd 2.37fF $ **FLOATING
C603 a_1026_45630.n176 gnd 6.33fF $ **FLOATING
C604 a_1026_45630.t10 gnd 2.37fF $ **FLOATING
C605 a_1026_45630.n177 gnd 6.33fF $ **FLOATING
C606 a_1026_45630.t140 gnd 2.37fF $ **FLOATING
C607 a_1026_45630.n178 gnd 6.33fF $ **FLOATING
C608 a_1026_45630.t97 gnd 2.37fF $ **FLOATING
C609 a_1026_45630.n179 gnd 3.52fF $ **FLOATING
C610 a_1026_45630.t27 gnd 2.37fF $ **FLOATING
C611 a_1026_45630.n180 gnd 2.94fF $ **FLOATING
C612 a_1026_45630.t65 gnd 6.88fF $ **FLOATING
C613 a_1026_45630.n181 gnd 8.73fF $ **FLOATING
C614 a_1026_45630.t198 gnd 2.37fF $ **FLOATING
C615 a_1026_45630.n182 gnd 6.45fF $ **FLOATING
C616 a_1026_45630.t92 gnd 2.37fF $ **FLOATING
C617 a_1026_45630.n183 gnd 6.33fF $ **FLOATING
C618 a_1026_45630.t39 gnd 2.37fF $ **FLOATING
C619 a_1026_45630.n184 gnd 6.33fF $ **FLOATING
C620 a_1026_45630.t175 gnd 2.37fF $ **FLOATING
C621 a_1026_45630.n185 gnd 6.33fF $ **FLOATING
C622 a_1026_45630.t22 gnd 2.37fF $ **FLOATING
C623 a_1026_45630.n186 gnd 6.33fF $ **FLOATING
C624 a_1026_45630.t168 gnd 2.37fF $ **FLOATING
C625 a_1026_45630.n187 gnd 6.33fF $ **FLOATING
C626 a_1026_45630.t103 gnd 2.37fF $ **FLOATING
C627 a_1026_45630.n188 gnd 6.33fF $ **FLOATING
C628 a_1026_45630.t53 gnd 2.37fF $ **FLOATING
C629 a_1026_45630.n189 gnd 3.52fF $ **FLOATING
C630 a_1026_45630.t186 gnd 2.37fF $ **FLOATING
C631 a_1026_45630.n190 gnd 2.93fF $ **FLOATING
C632 a_1026_45630.t66 gnd 6.91fF $ **FLOATING
C633 a_1026_45630.n191 gnd 8.75fF $ **FLOATING
C634 a_1026_45630.t199 gnd 2.37fF $ **FLOATING
C635 a_1026_45630.n192 gnd 6.45fF $ **FLOATING
C636 a_1026_45630.t93 gnd 2.37fF $ **FLOATING
C637 a_1026_45630.n193 gnd 6.33fF $ **FLOATING
C638 a_1026_45630.t40 gnd 2.37fF $ **FLOATING
C639 a_1026_45630.n194 gnd 6.33fF $ **FLOATING
C640 a_1026_45630.t176 gnd 2.37fF $ **FLOATING
C641 a_1026_45630.n195 gnd 6.33fF $ **FLOATING
C642 a_1026_45630.t23 gnd 2.37fF $ **FLOATING
C643 a_1026_45630.n196 gnd 6.33fF $ **FLOATING
C644 a_1026_45630.t169 gnd 2.37fF $ **FLOATING
C645 a_1026_45630.n197 gnd 6.33fF $ **FLOATING
C646 a_1026_45630.t104 gnd 2.37fF $ **FLOATING
C647 a_1026_45630.n198 gnd 6.33fF $ **FLOATING
C648 a_1026_45630.t54 gnd 2.37fF $ **FLOATING
C649 a_1026_45630.n199 gnd 3.52fF $ **FLOATING
C650 a_1026_45630.t187 gnd 2.37fF $ **FLOATING
C651 a_1026_45630.n200 gnd 3.08fF $ **FLOATING
C652 a_26690_784.n0 gnd 3.33fF $ **FLOATING
C653 a_23414_5032.t14 gnd 23.50fF $ **FLOATING
C654 a_23414_5032.t2 gnd 14.47fF $ **FLOATING
C655 a_26368_16652.t24 gnd 32.80fF $ **FLOATING
C656 a_26368_16652.n0 gnd 4.09fF $ **FLOATING
C657 Fvco_By4_QPH_bar.n0 gnd 21.37fF $ **FLOATING
C658 Fvco_By4_QPH_bar.n2 gnd 3.86fF $ **FLOATING
C659 Fvco_By4_QPH_bar.n3 gnd 3.48fF $ **FLOATING
C660 Fvco_By4_QPH_bar.n5 gnd 7.86fF $ **FLOATING
C661 a_34044_31208.n2 gnd 3.01fF $ **FLOATING
C662 a_34044_31208.n3 gnd 3.24fF $ **FLOATING
C663 a_34044_31208.t93 gnd 2.36fF $ **FLOATING
C664 a_34044_31208.n4 gnd 6.28fF $ **FLOATING
C665 a_34044_31208.t157 gnd 2.36fF $ **FLOATING
C666 a_34044_31208.n5 gnd 6.28fF $ **FLOATING
C667 a_34044_31208.t5 gnd 2.36fF $ **FLOATING
C668 a_34044_31208.n6 gnd 6.28fF $ **FLOATING
C669 a_34044_31208.t72 gnd 2.36fF $ **FLOATING
C670 a_34044_31208.n7 gnd 3.68fF $ **FLOATING
C671 a_34044_31208.t123 gnd 2.36fF $ **FLOATING
C672 a_34044_31208.n8 gnd 4.33fF $ **FLOATING
C673 a_34044_31208.n9 gnd 5.58fF $ **FLOATING
C674 a_34044_31208.t77 gnd 2.36fF $ **FLOATING
C675 a_34044_31208.n10 gnd 3.68fF $ **FLOATING
C676 a_34044_31208.t142 gnd 2.36fF $ **FLOATING
C677 a_34044_31208.n11 gnd 6.40fF $ **FLOATING
C678 a_34044_31208.t188 gnd 2.36fF $ **FLOATING
C679 a_34044_31208.n12 gnd 8.65fF $ **FLOATING
C680 a_34044_31208.t102 gnd 2.36fF $ **FLOATING
C681 a_34044_31208.t168 gnd 6.85fF $ **FLOATING
C682 a_34044_31208.t76 gnd 6.79fF $ **FLOATING
C683 a_34044_31208.n15 gnd 8.68fF $ **FLOATING
C684 a_34044_31208.t8 gnd 2.36fF $ **FLOATING
C685 a_34044_31208.n16 gnd 6.43fF $ **FLOATING
C686 a_34044_31208.t51 gnd 2.36fF $ **FLOATING
C687 a_34044_31208.n17 gnd 6.32fF $ **FLOATING
C688 a_34044_31208.t200 gnd 2.36fF $ **FLOATING
C689 a_34044_31208.n18 gnd 6.32fF $ **FLOATING
C690 a_34044_31208.t135 gnd 2.36fF $ **FLOATING
C691 a_34044_31208.n19 gnd 6.32fF $ **FLOATING
C692 a_34044_31208.t179 gnd 2.36fF $ **FLOATING
C693 a_34044_31208.n20 gnd 6.32fF $ **FLOATING
C694 a_34044_31208.t132 gnd 2.36fF $ **FLOATING
C695 a_34044_31208.n21 gnd 6.32fF $ **FLOATING
C696 a_34044_31208.t65 gnd 2.36fF $ **FLOATING
C697 a_34044_31208.n22 gnd 6.32fF $ **FLOATING
C698 a_34044_31208.t19 gnd 2.36fF $ **FLOATING
C699 a_34044_31208.n23 gnd 6.31fF $ **FLOATING
C700 a_34044_31208.t148 gnd 2.36fF $ **FLOATING
C701 a_34044_31208.n24 gnd 3.42fF $ **FLOATING
C702 a_34044_31208.t114 gnd 6.86fF $ **FLOATING
C703 a_34044_31208.n25 gnd 8.71fF $ **FLOATING
C704 a_34044_31208.t46 gnd 2.36fF $ **FLOATING
C705 a_34044_31208.n26 gnd 6.43fF $ **FLOATING
C706 a_34044_31208.t134 gnd 2.36fF $ **FLOATING
C707 a_34044_31208.n27 gnd 6.32fF $ **FLOATING
C708 a_34044_31208.t89 gnd 2.36fF $ **FLOATING
C709 a_34044_31208.n28 gnd 6.32fF $ **FLOATING
C710 a_34044_31208.t22 gnd 2.36fF $ **FLOATING
C711 a_34044_31208.n29 gnd 6.32fF $ **FLOATING
C712 a_34044_31208.t69 gnd 2.36fF $ **FLOATING
C713 a_34044_31208.n30 gnd 6.32fF $ **FLOATING
C714 a_34044_31208.t17 gnd 2.36fF $ **FLOATING
C715 a_34044_31208.n31 gnd 6.32fF $ **FLOATING
C716 a_34044_31208.t147 gnd 2.36fF $ **FLOATING
C717 a_34044_31208.n32 gnd 6.32fF $ **FLOATING
C718 a_34044_31208.t101 gnd 2.36fF $ **FLOATING
C719 a_34044_31208.n33 gnd 3.66fF $ **FLOATING
C720 a_34044_31208.t36 gnd 2.36fF $ **FLOATING
C721 a_34044_31208.n34 gnd 3.08fF $ **FLOATING
C722 a_34044_31208.t152 gnd 6.89fF $ **FLOATING
C723 a_34044_31208.n35 gnd 8.73fF $ **FLOATING
C724 a_34044_31208.t86 gnd 2.36fF $ **FLOATING
C725 a_34044_31208.n36 gnd 6.43fF $ **FLOATING
C726 a_34044_31208.t172 gnd 2.36fF $ **FLOATING
C727 a_34044_31208.n37 gnd 6.32fF $ **FLOATING
C728 a_34044_31208.t128 gnd 2.36fF $ **FLOATING
C729 a_34044_31208.n38 gnd 6.32fF $ **FLOATING
C730 a_34044_31208.t61 gnd 2.36fF $ **FLOATING
C731 a_34044_31208.n39 gnd 6.32fF $ **FLOATING
C732 a_34044_31208.t105 gnd 2.36fF $ **FLOATING
C733 a_34044_31208.n40 gnd 6.32fF $ **FLOATING
C734 a_34044_31208.t57 gnd 2.36fF $ **FLOATING
C735 a_34044_31208.n41 gnd 6.32fF $ **FLOATING
C736 a_34044_31208.t185 gnd 2.36fF $ **FLOATING
C737 a_34044_31208.n42 gnd 6.32fF $ **FLOATING
C738 a_34044_31208.t140 gnd 2.36fF $ **FLOATING
C739 a_34044_31208.n43 gnd 3.66fF $ **FLOATING
C740 a_34044_31208.t74 gnd 2.36fF $ **FLOATING
C741 a_34044_31208.n44 gnd 3.09fF $ **FLOATING
C742 a_34044_31208.t62 gnd 6.82fF $ **FLOATING
C743 a_34044_31208.n45 gnd 8.69fF $ **FLOATING
C744 a_34044_31208.t192 gnd 2.36fF $ **FLOATING
C745 a_34044_31208.n46 gnd 6.43fF $ **FLOATING
C746 a_34044_31208.t82 gnd 2.36fF $ **FLOATING
C747 a_34044_31208.n47 gnd 6.32fF $ **FLOATING
C748 a_34044_31208.t37 gnd 2.36fF $ **FLOATING
C749 a_34044_31208.n48 gnd 6.32fF $ **FLOATING
C750 a_34044_31208.t165 gnd 2.36fF $ **FLOATING
C751 a_34044_31208.n49 gnd 6.32fF $ **FLOATING
C752 a_34044_31208.t15 gnd 2.36fF $ **FLOATING
C753 a_34044_31208.n50 gnd 6.32fF $ **FLOATING
C754 a_34044_31208.t161 gnd 2.36fF $ **FLOATING
C755 a_34044_31208.n51 gnd 6.32fF $ **FLOATING
C756 a_34044_31208.t97 gnd 2.36fF $ **FLOATING
C757 a_34044_31208.n52 gnd 6.32fF $ **FLOATING
C758 a_34044_31208.t53 gnd 2.36fF $ **FLOATING
C759 a_34044_31208.n53 gnd 3.66fF $ **FLOATING
C760 a_34044_31208.t182 gnd 2.36fF $ **FLOATING
C761 a_34044_31208.n54 gnd 3.09fF $ **FLOATING
C762 a_34044_31208.t191 gnd 6.82fF $ **FLOATING
C763 a_34044_31208.n55 gnd 8.69fF $ **FLOATING
C764 a_34044_31208.t124 gnd 2.36fF $ **FLOATING
C765 a_34044_31208.n56 gnd 6.43fF $ **FLOATING
C766 a_34044_31208.t13 gnd 2.36fF $ **FLOATING
C767 a_34044_31208.n57 gnd 6.32fF $ **FLOATING
C768 a_34044_31208.t164 gnd 2.36fF $ **FLOATING
C769 a_34044_31208.n58 gnd 6.32fF $ **FLOATING
C770 a_34044_31208.t99 gnd 2.36fF $ **FLOATING
C771 a_34044_31208.n59 gnd 6.32fF $ **FLOATING
C772 a_34044_31208.t144 gnd 2.36fF $ **FLOATING
C773 a_34044_31208.n60 gnd 6.32fF $ **FLOATING
C774 a_34044_31208.t96 gnd 2.36fF $ **FLOATING
C775 a_34044_31208.n61 gnd 6.32fF $ **FLOATING
C776 a_34044_31208.t30 gnd 2.36fF $ **FLOATING
C777 a_34044_31208.n62 gnd 6.32fF $ **FLOATING
C778 a_34044_31208.t181 gnd 2.36fF $ **FLOATING
C779 a_34044_31208.n63 gnd 3.66fF $ **FLOATING
C780 a_34044_31208.t116 gnd 2.36fF $ **FLOATING
C781 a_34044_31208.n64 gnd 3.08fF $ **FLOATING
C782 a_34044_31208.t33 gnd 6.82fF $ **FLOATING
C783 a_34044_31208.n65 gnd 8.69fF $ **FLOATING
C784 a_34044_31208.t163 gnd 2.36fF $ **FLOATING
C785 a_34044_31208.n66 gnd 6.43fF $ **FLOATING
C786 a_34044_31208.t71 gnd 2.36fF $ **FLOATING
C787 a_34044_31208.n67 gnd 6.32fF $ **FLOATING
C788 a_34044_31208.t27 gnd 2.36fF $ **FLOATING
C789 a_34044_31208.n68 gnd 6.32fF $ **FLOATING
C790 a_34044_31208.t155 gnd 2.36fF $ **FLOATING
C791 a_34044_31208.n69 gnd 6.32fF $ **FLOATING
C792 a_34044_31208.t4 gnd 2.36fF $ **FLOATING
C793 a_34044_31208.n70 gnd 6.32fF $ **FLOATING
C794 a_34044_31208.t153 gnd 2.36fF $ **FLOATING
C795 a_34044_31208.n71 gnd 6.32fF $ **FLOATING
C796 a_34044_31208.t88 gnd 2.36fF $ **FLOATING
C797 a_34044_31208.n72 gnd 6.32fF $ **FLOATING
C798 a_34044_31208.t41 gnd 2.36fF $ **FLOATING
C799 a_34044_31208.n73 gnd 3.66fF $ **FLOATING
C800 a_34044_31208.t171 gnd 2.36fF $ **FLOATING
C801 a_34044_31208.n74 gnd 3.08fF $ **FLOATING
C802 a_34044_31208.t91 gnd 6.82fF $ **FLOATING
C803 a_34044_31208.n75 gnd 8.69fF $ **FLOATING
C804 a_34044_31208.t25 gnd 2.36fF $ **FLOATING
C805 a_34044_31208.n76 gnd 6.43fF $ **FLOATING
C806 a_34044_31208.t112 gnd 2.36fF $ **FLOATING
C807 a_34044_31208.n77 gnd 6.32fF $ **FLOATING
C808 a_34044_31208.t67 gnd 2.36fF $ **FLOATING
C809 a_34044_31208.n78 gnd 6.32fF $ **FLOATING
C810 a_34044_31208.t199 gnd 2.36fF $ **FLOATING
C811 a_34044_31208.n79 gnd 6.32fF $ **FLOATING
C812 a_34044_31208.t47 gnd 2.36fF $ **FLOATING
C813 a_34044_31208.n80 gnd 6.32fF $ **FLOATING
C814 a_34044_31208.t196 gnd 2.36fF $ **FLOATING
C815 a_34044_31208.n81 gnd 6.32fF $ **FLOATING
C816 a_34044_31208.t127 gnd 2.36fF $ **FLOATING
C817 a_34044_31208.n82 gnd 6.32fF $ **FLOATING
C818 a_34044_31208.t81 gnd 2.36fF $ **FLOATING
C819 a_34044_31208.n83 gnd 3.66fF $ **FLOATING
C820 a_34044_31208.t12 gnd 2.36fF $ **FLOATING
C821 a_34044_31208.n84 gnd 3.08fF $ **FLOATING
C822 a_34044_31208.t109 gnd 6.86fF $ **FLOATING
C823 a_34044_31208.n85 gnd 8.71fF $ **FLOATING
C824 a_34044_31208.t42 gnd 2.36fF $ **FLOATING
C825 a_34044_31208.n86 gnd 6.43fF $ **FLOATING
C826 a_34044_31208.t131 gnd 2.36fF $ **FLOATING
C827 a_34044_31208.n87 gnd 6.32fF $ **FLOATING
C828 a_34044_31208.t84 gnd 2.36fF $ **FLOATING
C829 a_34044_31208.n88 gnd 6.32fF $ **FLOATING
C830 a_34044_31208.t18 gnd 2.36fF $ **FLOATING
C831 a_34044_31208.n89 gnd 6.32fF $ **FLOATING
C832 a_34044_31208.t66 gnd 2.36fF $ **FLOATING
C833 a_34044_31208.n90 gnd 6.32fF $ **FLOATING
C834 a_34044_31208.t11 gnd 2.36fF $ **FLOATING
C835 a_34044_31208.n91 gnd 6.32fF $ **FLOATING
C836 a_34044_31208.t141 gnd 2.36fF $ **FLOATING
C837 a_34044_31208.n92 gnd 6.32fF $ **FLOATING
C838 a_34044_31208.t98 gnd 2.36fF $ **FLOATING
C839 a_34044_31208.n93 gnd 3.66fF $ **FLOATING
C840 a_34044_31208.t31 gnd 2.36fF $ **FLOATING
C841 a_34044_31208.n94 gnd 3.08fF $ **FLOATING
C842 a_34044_31208.t20 gnd 6.82fF $ **FLOATING
C843 a_34044_31208.n95 gnd 8.69fF $ **FLOATING
C844 a_34044_31208.t149 gnd 2.36fF $ **FLOATING
C845 a_34044_31208.n96 gnd 6.43fF $ **FLOATING
C846 a_34044_31208.t39 gnd 2.36fF $ **FLOATING
C847 a_34044_31208.n97 gnd 6.32fF $ **FLOATING
C848 a_34044_31208.t190 gnd 2.36fF $ **FLOATING
C849 a_34044_31208.n98 gnd 6.32fF $ **FLOATING
C850 a_34044_31208.t122 gnd 2.36fF $ **FLOATING
C851 a_34044_31208.n99 gnd 6.32fF $ **FLOATING
C852 a_34044_31208.t169 gnd 2.36fF $ **FLOATING
C853 a_34044_31208.n100 gnd 6.32fF $ **FLOATING
C854 a_34044_31208.t118 gnd 2.36fF $ **FLOATING
C855 a_34044_31208.n101 gnd 6.32fF $ **FLOATING
C856 a_34044_31208.t54 gnd 2.36fF $ **FLOATING
C857 a_34044_31208.n102 gnd 6.32fF $ **FLOATING
C858 a_34044_31208.t6 gnd 2.36fF $ **FLOATING
C859 a_34044_31208.n103 gnd 3.66fF $ **FLOATING
C860 a_34044_31208.t138 gnd 2.36fF $ **FLOATING
C861 a_34044_31208.n104 gnd 3.09fF $ **FLOATING
C862 a_34044_31208.t59 gnd 6.86fF $ **FLOATING
C863 a_34044_31208.n105 gnd 8.71fF $ **FLOATING
C864 a_34044_31208.t187 gnd 2.36fF $ **FLOATING
C865 a_34044_31208.n106 gnd 6.43fF $ **FLOATING
C866 a_34044_31208.t79 gnd 2.36fF $ **FLOATING
C867 a_34044_31208.n107 gnd 6.32fF $ **FLOATING
C868 a_34044_31208.t32 gnd 2.36fF $ **FLOATING
C869 a_34044_31208.n108 gnd 6.32fF $ **FLOATING
C870 a_34044_31208.t162 gnd 2.36fF $ **FLOATING
C871 a_34044_31208.n109 gnd 6.32fF $ **FLOATING
C872 a_34044_31208.t10 gnd 2.36fF $ **FLOATING
C873 a_34044_31208.n110 gnd 6.32fF $ **FLOATING
C874 a_34044_31208.t158 gnd 2.36fF $ **FLOATING
C875 a_34044_31208.n111 gnd 6.32fF $ **FLOATING
C876 a_34044_31208.t94 gnd 2.36fF $ **FLOATING
C877 a_34044_31208.n112 gnd 6.32fF $ **FLOATING
C878 a_34044_31208.t49 gnd 2.36fF $ **FLOATING
C879 a_34044_31208.n113 gnd 3.66fF $ **FLOATING
C880 a_34044_31208.t177 gnd 2.36fF $ **FLOATING
C881 a_34044_31208.n114 gnd 3.08fF $ **FLOATING
C882 a_34044_31208.t58 gnd 6.82fF $ **FLOATING
C883 a_34044_31208.n115 gnd 8.69fF $ **FLOATING
C884 a_34044_31208.t186 gnd 2.36fF $ **FLOATING
C885 a_34044_31208.n116 gnd 6.43fF $ **FLOATING
C886 a_34044_31208.t29 gnd 2.36fF $ **FLOATING
C887 a_34044_31208.n117 gnd 6.32fF $ **FLOATING
C888 a_34044_31208.t180 gnd 2.36fF $ **FLOATING
C889 a_34044_31208.n118 gnd 6.32fF $ **FLOATING
C890 a_34044_31208.t115 gnd 2.36fF $ **FLOATING
C891 a_34044_31208.n119 gnd 6.32fF $ **FLOATING
C892 a_34044_31208.t159 gnd 2.36fF $ **FLOATING
C893 a_34044_31208.n120 gnd 6.32fF $ **FLOATING
C894 a_34044_31208.t110 gnd 2.36fF $ **FLOATING
C895 a_34044_31208.n121 gnd 6.32fF $ **FLOATING
C896 a_34044_31208.t44 gnd 2.36fF $ **FLOATING
C897 a_34044_31208.n122 gnd 6.32fF $ **FLOATING
C898 a_34044_31208.t198 gnd 2.36fF $ **FLOATING
C899 a_34044_31208.n123 gnd 3.66fF $ **FLOATING
C900 a_34044_31208.t130 gnd 2.36fF $ **FLOATING
C901 a_34044_31208.n124 gnd 3.08fF $ **FLOATING
C902 a_34044_31208.t50 gnd 6.86fF $ **FLOATING
C903 a_34044_31208.n125 gnd 8.71fF $ **FLOATING
C904 a_34044_31208.t178 gnd 2.36fF $ **FLOATING
C905 a_34044_31208.n126 gnd 6.43fF $ **FLOATING
C906 a_34044_31208.t70 gnd 2.36fF $ **FLOATING
C907 a_34044_31208.n127 gnd 6.32fF $ **FLOATING
C908 a_34044_31208.t24 gnd 2.36fF $ **FLOATING
C909 a_34044_31208.n128 gnd 6.32fF $ **FLOATING
C910 a_34044_31208.t154 gnd 2.36fF $ **FLOATING
C911 a_34044_31208.n129 gnd 6.32fF $ **FLOATING
C912 a_34044_31208.t201 gnd 2.36fF $ **FLOATING
C913 a_34044_31208.n130 gnd 6.32fF $ **FLOATING
C914 a_34044_31208.t150 gnd 2.36fF $ **FLOATING
C915 a_34044_31208.n131 gnd 6.32fF $ **FLOATING
C916 a_34044_31208.t83 gnd 2.36fF $ **FLOATING
C917 a_34044_31208.n132 gnd 6.32fF $ **FLOATING
C918 a_34044_31208.t38 gnd 2.36fF $ **FLOATING
C919 a_34044_31208.n133 gnd 3.66fF $ **FLOATING
C920 a_34044_31208.t167 gnd 2.36fF $ **FLOATING
C921 a_34044_31208.n134 gnd 3.08fF $ **FLOATING
C922 a_34044_31208.t90 gnd 6.82fF $ **FLOATING
C923 a_34044_31208.n135 gnd 8.69fF $ **FLOATING
C924 a_34044_31208.t23 gnd 2.36fF $ **FLOATING
C925 a_34044_31208.n136 gnd 6.43fF $ **FLOATING
C926 a_34044_31208.t108 gnd 2.36fF $ **FLOATING
C927 a_34044_31208.n137 gnd 6.32fF $ **FLOATING
C928 a_34044_31208.t64 gnd 2.36fF $ **FLOATING
C929 a_34044_31208.n138 gnd 6.32fF $ **FLOATING
C930 a_34044_31208.t197 gnd 2.36fF $ **FLOATING
C931 a_34044_31208.n139 gnd 6.32fF $ **FLOATING
C932 a_34044_31208.t43 gnd 2.36fF $ **FLOATING
C933 a_34044_31208.n140 gnd 6.32fF $ **FLOATING
C934 a_34044_31208.t189 gnd 2.36fF $ **FLOATING
C935 a_34044_31208.n141 gnd 6.32fF $ **FLOATING
C936 a_34044_31208.t121 gnd 2.36fF $ **FLOATING
C937 a_34044_31208.n142 gnd 6.32fF $ **FLOATING
C938 a_34044_31208.t78 gnd 2.36fF $ **FLOATING
C939 a_34044_31208.n143 gnd 3.66fF $ **FLOATING
C940 a_34044_31208.t9 gnd 2.36fF $ **FLOATING
C941 a_34044_31208.n144 gnd 3.09fF $ **FLOATING
C942 a_34044_31208.t173 gnd 6.80fF $ **FLOATING
C943 a_34044_31208.n145 gnd 8.68fF $ **FLOATING
C944 a_34044_31208.t103 gnd 2.36fF $ **FLOATING
C945 a_34044_31208.n146 gnd 6.43fF $ **FLOATING
C946 a_34044_31208.t195 gnd 2.36fF $ **FLOATING
C947 a_34044_31208.n147 gnd 6.32fF $ **FLOATING
C948 a_34044_31208.t146 gnd 2.36fF $ **FLOATING
C949 a_34044_31208.n148 gnd 6.32fF $ **FLOATING
C950 a_34044_31208.t80 gnd 2.36fF $ **FLOATING
C951 a_34044_31208.n149 gnd 6.32fF $ **FLOATING
C952 a_34044_31208.t129 gnd 2.36fF $ **FLOATING
C953 a_34044_31208.n150 gnd 6.32fF $ **FLOATING
C954 a_34044_31208.t75 gnd 2.36fF $ **FLOATING
C955 a_34044_31208.n151 gnd 6.32fF $ **FLOATING
C956 a_34044_31208.t7 gnd 2.36fF $ **FLOATING
C957 a_34044_31208.n152 gnd 6.32fF $ **FLOATING
C958 a_34044_31208.t160 gnd 2.36fF $ **FLOATING
C959 a_34044_31208.n153 gnd 3.66fF $ **FLOATING
C960 a_34044_31208.t95 gnd 2.36fF $ **FLOATING
C961 a_34044_31208.n154 gnd 3.08fF $ **FLOATING
C962 a_34044_31208.t14 gnd 6.86fF $ **FLOATING
C963 a_34044_31208.n155 gnd 8.71fF $ **FLOATING
C964 a_34044_31208.t143 gnd 2.36fF $ **FLOATING
C965 a_34044_31208.n156 gnd 6.43fF $ **FLOATING
C966 a_34044_31208.t35 gnd 2.36fF $ **FLOATING
C967 a_34044_31208.n157 gnd 6.32fF $ **FLOATING
C968 a_34044_31208.t184 gnd 2.36fF $ **FLOATING
C969 a_34044_31208.n158 gnd 6.32fF $ **FLOATING
C970 a_34044_31208.t119 gnd 2.36fF $ **FLOATING
C971 a_34044_31208.n159 gnd 6.32fF $ **FLOATING
C972 a_34044_31208.t166 gnd 2.36fF $ **FLOATING
C973 a_34044_31208.n160 gnd 6.32fF $ **FLOATING
C974 a_34044_31208.t117 gnd 2.36fF $ **FLOATING
C975 a_34044_31208.n161 gnd 6.32fF $ **FLOATING
C976 a_34044_31208.t52 gnd 2.36fF $ **FLOATING
C977 a_34044_31208.n162 gnd 6.32fF $ **FLOATING
C978 a_34044_31208.t202 gnd 2.36fF $ **FLOATING
C979 a_34044_31208.n163 gnd 3.66fF $ **FLOATING
C980 a_34044_31208.t136 gnd 2.36fF $ **FLOATING
C981 a_34044_31208.n164 gnd 3.08fF $ **FLOATING
C982 a_34044_31208.t120 gnd 6.83fF $ **FLOATING
C983 a_34044_31208.n165 gnd 8.70fF $ **FLOATING
C984 a_34044_31208.t55 gnd 2.36fF $ **FLOATING
C985 a_34044_31208.n166 gnd 6.43fF $ **FLOATING
C986 a_34044_31208.t92 gnd 2.36fF $ **FLOATING
C987 a_34044_31208.n167 gnd 6.32fF $ **FLOATING
C988 a_34044_31208.t48 gnd 2.36fF $ **FLOATING
C989 a_34044_31208.n168 gnd 6.32fF $ **FLOATING
C990 a_34044_31208.t176 gnd 2.36fF $ **FLOATING
C991 a_34044_31208.n169 gnd 6.32fF $ **FLOATING
C992 a_34044_31208.t28 gnd 2.36fF $ **FLOATING
C993 a_34044_31208.n170 gnd 6.32fF $ **FLOATING
C994 a_34044_31208.t174 gnd 2.36fF $ **FLOATING
C995 a_34044_31208.n171 gnd 6.32fF $ **FLOATING
C996 a_34044_31208.t107 gnd 2.36fF $ **FLOATING
C997 a_34044_31208.n172 gnd 6.32fF $ **FLOATING
C998 a_34044_31208.t63 gnd 2.36fF $ **FLOATING
C999 a_34044_31208.n173 gnd 3.66fF $ **FLOATING
C1000 a_34044_31208.t194 gnd 2.36fF $ **FLOATING
C1001 a_34044_31208.n174 gnd 3.08fF $ **FLOATING
C1002 a_34044_31208.t203 gnd 6.86fF $ **FLOATING
C1003 a_34044_31208.n175 gnd 8.71fF $ **FLOATING
C1004 a_34044_31208.t137 gnd 2.36fF $ **FLOATING
C1005 a_34044_31208.n176 gnd 6.43fF $ **FLOATING
C1006 a_34044_31208.t26 gnd 2.36fF $ **FLOATING
C1007 a_34044_31208.n177 gnd 6.32fF $ **FLOATING
C1008 a_34044_31208.t175 gnd 2.36fF $ **FLOATING
C1009 a_34044_31208.n178 gnd 6.32fF $ **FLOATING
C1010 a_34044_31208.t111 gnd 2.36fF $ **FLOATING
C1011 a_34044_31208.n179 gnd 6.32fF $ **FLOATING
C1012 a_34044_31208.t156 gnd 2.36fF $ **FLOATING
C1013 a_34044_31208.n180 gnd 6.32fF $ **FLOATING
C1014 a_34044_31208.t106 gnd 2.36fF $ **FLOATING
C1015 a_34044_31208.n181 gnd 6.32fF $ **FLOATING
C1016 a_34044_31208.t40 gnd 2.36fF $ **FLOATING
C1017 a_34044_31208.n182 gnd 6.32fF $ **FLOATING
C1018 a_34044_31208.t193 gnd 2.36fF $ **FLOATING
C1019 a_34044_31208.n183 gnd 3.66fF $ **FLOATING
C1020 a_34044_31208.t125 gnd 2.36fF $ **FLOATING
C1021 a_34044_31208.n184 gnd 3.09fF $ **FLOATING
C1022 a_34044_31208.t113 gnd 6.86fF $ **FLOATING
C1023 a_34044_31208.n185 gnd 8.71fF $ **FLOATING
C1024 a_34044_31208.t45 gnd 2.36fF $ **FLOATING
C1025 a_34044_31208.n186 gnd 6.43fF $ **FLOATING
C1026 a_34044_31208.t133 gnd 2.36fF $ **FLOATING
C1027 a_34044_31208.n187 gnd 6.32fF $ **FLOATING
C1028 a_34044_31208.t87 gnd 2.36fF $ **FLOATING
C1029 a_34044_31208.n188 gnd 6.32fF $ **FLOATING
C1030 a_34044_31208.t21 gnd 2.36fF $ **FLOATING
C1031 a_34044_31208.n189 gnd 6.32fF $ **FLOATING
C1032 a_34044_31208.t68 gnd 2.36fF $ **FLOATING
C1033 a_34044_31208.n190 gnd 6.32fF $ **FLOATING
C1034 a_34044_31208.t16 gnd 2.36fF $ **FLOATING
C1035 a_34044_31208.n191 gnd 6.32fF $ **FLOATING
C1036 a_34044_31208.t145 gnd 2.36fF $ **FLOATING
C1037 a_34044_31208.n192 gnd 6.32fF $ **FLOATING
C1038 a_34044_31208.t100 gnd 2.36fF $ **FLOATING
C1039 a_34044_31208.n193 gnd 3.66fF $ **FLOATING
C1040 a_34044_31208.t34 gnd 2.36fF $ **FLOATING
C1041 a_34044_31208.n194 gnd 3.08fF $ **FLOATING
C1042 a_34044_31208.t151 gnd 6.86fF $ **FLOATING
C1043 a_34044_31208.n195 gnd 8.71fF $ **FLOATING
C1044 a_34044_31208.t85 gnd 2.36fF $ **FLOATING
C1045 a_34044_31208.n196 gnd 6.43fF $ **FLOATING
C1046 a_34044_31208.t170 gnd 2.36fF $ **FLOATING
C1047 a_34044_31208.n197 gnd 6.32fF $ **FLOATING
C1048 a_34044_31208.t126 gnd 2.36fF $ **FLOATING
C1049 a_34044_31208.n198 gnd 6.32fF $ **FLOATING
C1050 a_34044_31208.t60 gnd 2.36fF $ **FLOATING
C1051 a_34044_31208.n199 gnd 6.32fF $ **FLOATING
C1052 a_34044_31208.t104 gnd 2.36fF $ **FLOATING
C1053 a_34044_31208.n200 gnd 6.32fF $ **FLOATING
C1054 a_34044_31208.t56 gnd 2.36fF $ **FLOATING
C1055 a_34044_31208.n201 gnd 6.32fF $ **FLOATING
C1056 a_34044_31208.t183 gnd 2.36fF $ **FLOATING
C1057 a_34044_31208.n202 gnd 6.32fF $ **FLOATING
C1058 a_34044_31208.t139 gnd 2.36fF $ **FLOATING
C1059 a_34044_31208.n203 gnd 3.66fF $ **FLOATING
C1060 a_34044_31208.t73 gnd 2.36fF $ **FLOATING
