* NGSPICE file created from loopwithesd.ext - technology: sky130A

X0 Fvco_By4_QPH_bar.t1 a_66167_26022# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X1 a_28994_17218# a_26368_16652.t2 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X2 a_26690_784.t1 a_23414_5032.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X3 vdd Vso1b a_4226_11420# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X4 vinit.t39 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X5 gnd gnd vinit.t19 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X6 a_28220_17218# a_26368_16652.t3 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X7 a_29510_17218# a_26368_16652.t4 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X8 a_23403_5596# a_14188_14050.t2 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X9 a_22629_5596# a_14188_14050.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X10 a_49874_4150.t1 a_49874_4150.t0 a_54950_4814# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.856e+11p ps=1.57e+06u w=1.28e+06u l=8e+06u
X11 a_50320_14126# Fvco_By4_QPH.t2 a_55602_11692# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=1.98421e+11p ps=1.49053e+06u w=1e+06u l=150000u
X12 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X13 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X14 a_29510_17218# a_26368_16652.t5 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X15 a_28994_5597# a_26036_4988.t2 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X16 a_22887_5596# a_14188_14050.t4 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X17 a_54950_4814# a_49874_4150.t4 a_53292_4814# gnd sky130_fd_pr__nfet_01v8 ad=1.856e+11p pd=1.57e+06u as=1.856e+11p ps=1.57e+06u w=1.28e+06u l=8e+06u
X18 a_26847_11500# a_25099_11445.t2 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X19 vdd a_66167_26022# a_66154_26414# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X20 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X21 a_24177_5596# a_14188_14050.t5 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X22 gnd a_17685_3840.t17 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X23 a_22629_11500# a_14266_8900.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X24 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X25 gnd a_17685_3840.t18 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X26 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X27 a_66357_25280# RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=6.405e+10p pd=725000u as=9.2007e+10p ps=682276u w=420000u l=150000u
X28 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X29 vdd a_63529_26290# a_63419_26414# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=1.134e+11p ps=1.1e+06u w=420000u l=150000u
X30 a_28736_5597# a_26036_4988.t3 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X31 a_77268_24654# a_77242_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X32 a_26847_11500# a_25099_11445.t3 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X33 a_29510_5597# a_26036_4988.t4 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X34 gnd Vso3b a_8744_13422# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X35 gnd a_17685_3840.t19 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X36 gnd Vso5b a_8748_12270# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X37 a_26847_11500# a_25099_11445.t4 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X38 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X39 a_23919_5596# a_14188_14050.t6 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X40 a_28994_5597# a_26036_4988.t5 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X41 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X42 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X43 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X44 a_52052_20860.t18 a_56334_20860.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X45 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X46 a_26847_11500# a_25099_11445.t5 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X47 a_23156_5032.t7 a_14188_14050.t7 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X48 vbiasr.t40 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X49 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X50 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X51 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X52 a_28736_17218# a_26368_16652.t6 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X53 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X54 a_65546_25646# RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=9.08803e+10p ps=655615u w=420000u l=150000u
X55 a_25299_17217# a_23436_16644.t2 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X56 a_26847_17217# a_23436_16644.t3 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X57 a_28736_17218# a_26368_16652.t7 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X58 a_25815_5596# a_23414_5032.t3 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X59 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X60 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X61 a_51276_14152# Fvco_By4_QPH.t3 a_51636_13108# gnd sky130_fd_pr__nfet_01v8 ad=2.07143e+11p pd=1.67714e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X62 gnd a_17685_3840.t20 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X63 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X64 a_63311_26048# a_62795_26048# a_63216_26048# gnd sky130_fd_pr__nfet_01v8 ad=5.94e+10p pd=690000u as=6.09231e+10p ps=687692u w=360000u l=150000u
X65 a_23145_5596# a_14188_14050.t8 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X66 vdd vdd vinit.t38 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X67 a_26331_11500# a_25099_11445.t6 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X68 a_28478_5597# a_26036_4988.t6 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X69 vbiasr.t39 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X70 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X71 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X72 a_29252_5597# a_26036_4988.t7 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X73 vdd CLK_IN a_4288_11534# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X74 a_25778_4988.t6 a_23414_5032.t4 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X75 a_26331_11500# a_25099_11445.t7 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X76 gnd a_17685_3840.t21 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X77 a_23145_17217# Fvco.t2 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X78 vinit.t18 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X79 a_28220_17218# a_26368_16652.t8 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X80 a_23145_17217# Fvco.t3 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X81 a_52052_20860.t8 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X82 a_56602_11692# vbiasob.t3 a_56272_15934.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=2e+06u
X83 a_27962_5597# a_26036_4988.t8 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X84 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X85 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X86 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X87 vbiasbuffer.t0 a_49874_4150.t5 a_54966_2992# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.9575e+11p ps=1.64e+06u w=1.35e+06u l=8e+06u
X88 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X89 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X90 a_26331_17217# a_23436_16644.t4 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X91 a_28220_17218# a_26368_16652.t9 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X92 vbiasob.t0 a_57726_5786.t5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.23446e+11p ps=1.65695e+06u w=1.02e+06u l=1e+06u
X93 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X94 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X95 a_25557_11500# a_25099_11445.t8 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X96 a_25557_5596# a_23414_5032.t5 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X97 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X98 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X99 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X100 a_22887_5596# a_14188_14050.t9 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X101 a_23661_5596# a_14188_14050.t10 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X102 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X103 a_26847_5596# a_23414_5032.t6 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X104 a_28578_5014.t6 a_26036_4988.t9 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X105 vctrl CLK_BY_4_IPH_BAR.t2 a_34590_30714# gnd sky130_fd_pr__nfet_01v8 ad=3.012e+11p pd=2.62e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X106 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X107 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X108 a_28220_5597# a_26036_4988.t10 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X109 gnd a_17685_3840.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X110 a_24177_11500# a_14266_8900.t3 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X111 a_50583_13108.t0 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X112 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X113 a_25557_11500# a_25099_11445.t9 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X114 a_52052_20860.t17 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X115 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X116 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X117 a_23403_5596# a_14188_14050.t11 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X118 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X119 a_29252_11501# a_27762_11446.t2 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X120 a_25557_11500# a_25099_11445.t10 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X121 a_25299_5596# a_23414_5032.t7 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X122 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X123 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X124 vdd vdd vinit.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X125 a_49932_4124.t2 a_49932_4124.t1 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=2e+07u
X126 a_28994_5597# a_26036_4988.t11 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X127 a_25557_11500# a_25099_11445.t11 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X128 vdd vdd vbiasr.t38 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X129 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X130 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X131 a_65438_25280# a_65088_25280# a_65343_25280# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.245e+10p pd=765000u as=6.51e+10p ps=730000u w=420000u l=150000u
X132 a_66346_26048# RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=6.405e+10p pd=725000u as=9.2007e+10p ps=682276u w=420000u l=150000u
X133 a_26589_5596# a_23414_5032.t8 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X134 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X135 a_65656_25522# a_65438_25280# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.722e+11p pd=1.58e+06u as=1.81761e+11p ps=1.31123e+06u w=840000u l=150000u
X136 a_24177_11500# a_14266_8900.t4 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X137 a_44752_16348.t2 a_51138_19904.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X138 a_25557_17217# a_23436_16644.t5 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X139 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X140 vinit.t17 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X141 a_24177_11500# a_14266_8900.t5 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X142 a_27962_11501# a_27762_11446.t3 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X143 vdd vdd vbiasr.t37 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X144 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X145 a_14832_12082.t1 a_14188_14050.t12 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X146 a_29252_11501# a_27762_11446.t4 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X147 a_56602_11692# a_51636_13108# a_52052_20860.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X148 a_29510_5597# a_26036_4988.t12 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X149 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X150 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X151 a_24177_11500# a_14266_8900.t6 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X152 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X153 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X154 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X155 a_66003_25280# a_64922_25280# a_65656_25522# vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=8.61e+10p ps=790000u w=420000u l=150000u
X156 a_29252_11501# a_27762_11446.t5 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X157 vdd a_56334_19906# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X158 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X159 a_26073_5596# a_23414_5032.t9 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X160 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X161 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X162 a_24177_17217# Fvco.t4 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X163 a_29252_11501# a_27762_11446.t6 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X164 a_26847_17217# a_23436_16644.t6 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X165 a_23160_10936.t6 a_14266_8900.t7 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X166 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X167 gnd Vso7b a_8748_11114# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X168 a_29252_17218# a_26368_16652.t10 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X169 a_23661_11500# a_14266_8900.t8 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X170 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X171 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X172 a_26847_17217# a_23436_16644.t7 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X173 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X174 a_23661_11500# a_14266_8900.t9 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X175 a_25815_5596# a_23414_5032.t10 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X176 a_23919_11500# a_14266_8900.t10 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X177 a_26331_5596# a_23414_5032.t11 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X178 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X179 a_77586_24654# a_77560_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X180 a_55602_11692# a_51041_13108# a_52052_20860.t16 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X181 a_42574_15624# Fvco_By4_QPH_bar.t2 a_42550_16062# vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X182 a_29252_5597# a_26036_4988.t13 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X183 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X184 a_53308_3580# a_49874_4150.t6 vbiasr.t20 gnd sky130_fd_pr__nfet_01v8 ad=7.0035e+11p pd=5.12e+06u as=0p ps=0u w=4.83e+06u l=8e+06u
X185 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X186 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X187 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X188 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X189 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X190 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X191 a_23661_17217# Fvco.t5 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X192 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X193 a_26331_17217# a_23436_16644.t8 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X194 a_22887_11500# a_14266_8900.t11 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X195 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X196 CLK_BY_4_IPH_BAR.t1 a_66742_25280# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X197 a_28438_10874.t6 a_27762_11446.t7 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X198 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X199 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X200 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X201 gnd a_17685_3840.t23 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X202 a_26331_17217# a_23436_16644.t9 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X203 a_23919_11500# a_14266_8900.t12 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X204 gnd gnd vbiasr.t19 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X205 gnd a_17685_3840.t24 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X206 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X207 a_28438_10874.t5 a_27762_11446.t8 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X208 a_25557_5596# a_23414_5032.t12 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X209 vinit.t36 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X210 a_23919_11500# a_14266_8900.t13 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X211 a_65438_25280# a_64922_25280# a_65343_25280# gnd sky130_fd_pr__nfet_01v8 ad=5.94e+10p pd=690000u as=6.09231e+10p ps=687692u w=360000u l=150000u
X212 a_23919_11500# a_14266_8900.t14 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X213 a_63573_26048# a_63529_26290# a_63407_26048# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.50877e+11p ps=1.18462e+06u w=420000u l=150000u
X214 gnd a_17685_3840.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X215 a_22887_11500# a_14266_8900.t15 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X216 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X217 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X218 a_14910_6932.t1 a_14266_8900.t16 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X219 a_28622_16652# a_26368_16652.t11 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X220 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X221 gnd Vso4b a_8740_12844# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X222 a_4314_11564# a_4288_11534# a_4314_11468# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X223 a_23919_17217# Fvco.t4 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X224 a_22887_11500# a_14266_8900.t17 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X225 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X226 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X227 gnd a_17685_3840.t26 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X228 gnd a_17685_3840.t27 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X229 vdd a_4288_11918# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X230 a_23403_11500# a_14266_8900.t18 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X231 a_22887_11500# a_14266_8900.t19 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X232 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X233 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X234 CLK_BY_2_BAR a_64615_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X235 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X236 a_23403_11500# a_14266_8900.t20 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X237 a_26016_10878.t6 a_25099_11445.t12 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X238 a_25299_5596# a_23414_5032.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X239 a_22887_17217# Fvco.t4 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X240 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X241 a_64725_25280# CLK_BY_2_BAR vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.35e+11p pd=1.27e+06u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X242 a_28622_16652# a_26368_16652.t12 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X243 a_25557_17217# a_23436_16644.t10 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X244 a_34590_30714# CLK_BY_4_IPH.t2 vctrl vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X245 gnd a_17685_3840.t28 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X246 a_25557_17217# a_23436_16644.t11 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X247 a_26073_11500# a_25099_11445.t13 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X248 gnd a_57726_5786.t2 a_57726_5786.t3 gnd sky130_fd_pr__nfet_01v8 ad=6.57193e+11p pd=4.8734e+06u as=0p ps=0u w=3e+06u l=1e+06u
X249 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X250 a_23403_17217# Fvco.t4 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X251 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X252 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X253 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X254 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X255 a_22629_11500# a_14266_8900.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X256 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X257 gnd gnd vbiasr.t18 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X258 a_49932_4124.t0 a_49874_4150.t7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.80402e+11p ps=2.07932e+06u w=1.28e+06u l=8e+06u
X259 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X260 a_24177_17217# Fvco.t6 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X261 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X262 a_24177_17217# Fvco.t7 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X263 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X264 gnd RESET a_63573_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=4.41e+10p ps=630000u w=420000u l=150000u
X265 a_29252_17218# a_26368_16652.t13 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X266 vbiasob.t2 vbiasob.t1 a_54448_7822.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X267 Vso1b a_24410_25128.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X268 a_28478_11501# a_27762_11446.t9 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X269 a_29252_17218# a_26368_16652.t14 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X270 a_22629_11500# a_14266_8900.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X271 a_23308_802.t0 Fvco.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X272 vbiasr.t17 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X273 a_26368_16652.t1 a_23436_16644.t12 a_26110_16652# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X274 a_28478_11501# a_27762_11446.t10 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X275 a_24177_5596# a_14188_14050.t13 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X276 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.19064e+11p pd=1.62447e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X277 vdd vdd vinit.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X278 a_22629_11500# a_14266_8900.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X279 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X280 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X281 a_77268_24654# a_77242_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X282 a_22629_11500# a_14266_8900.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X283 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X284 a_23661_17217# Fvco.t9 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X285 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X286 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X287 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X288 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X289 gnd Vso1b a_8744_9386# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X290 a_28478_17218# a_26368_16652.t15 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X291 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X292 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X293 a_22629_17217# Fvco.t4 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X294 a_23661_17217# Fvco.t10 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X295 a_26036_4988.t0 a_23414_5032.t14 a_17685_3840.t6 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X296 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X297 vdd a_4226_11420# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X298 gnd a_64725_25280# a_64922_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X299 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X300 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X301 vdd a_4226_12188# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X302 a_25815_11500# a_25099_11445.t14 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X303 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X304 gnd gnd vinit.t16 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X305 a_32948_24994.t1 a_27762_11446.t11 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X306 Vso2b a_28790_25040.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X307 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X308 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X309 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X310 a_28478_17218# a_26368_16652.t16 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X311 vbiasr.t16 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X312 a_28622_16652# a_26368_16652.t17 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X313 a_23145_5596# a_14188_14050.t14 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X314 a_23919_17217# Fvco.t11 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X315 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X316 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X317 gnd a_17685_3840.t29 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X318 a_28622_16652# a_26368_16652.t18 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X319 gnd gnd vinit.t15 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X320 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X321 vdd a_66167_26022# a_66731_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X322 a_23919_17217# Fvco.t12 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X323 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X324 a_14910_6932.t0 a_14266_8900.t25 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X325 gnd a_17685_3840.t30 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X326 a_52052_20860.t6 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X327 gnd a_17685_3840.t31 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X328 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X329 vbiasr.t15 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X330 a_51276_14152# a_51334_14126# z.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X331 vdd a_65992_26048# a_66167_26022# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X332 vdd Vso6b a_4226_11804# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X333 a_22887_17217# Fvco.t13 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X334 a_29510_11501# a_27762_11446.t12 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X335 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X336 a_27962_5597# a_26036_4988.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X337 a_22887_17217# Fvco.t14 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X338 a_51532_4150.t1 a_51532_4150.t0 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.59194e+11p ps=2.59124e+06u w=1.66e+06u l=4e+06u
X339 vdd a_65656_25522# a_65546_25646# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=1.134e+11p ps=1.1e+06u w=420000u l=150000u
X340 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X341 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X342 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X343 vdd CLK_BY_2_BAR a_64911_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X344 a_56602_11692# a_51636_13108# a_52052_20860.t5 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X345 vdd a_50032_16080.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X346 a_23403_17217# Fvco.t15 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X347 a_23661_5596# a_14188_14050.t15 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X348 a_22887_5596# a_14188_14050.t16 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X349 a_50511_16072.t5 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X350 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X351 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X352 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X353 a_64038_26414# a_62961_26048# a_63876_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=5.88e+10p ps=700000u w=420000u l=150000u
X354 a_23403_17217# Fvco.t16 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X355 a_23919_5596# a_14188_14050.t17 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X356 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X357 vdd a_51138_19904.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X358 z.t6 a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X359 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X360 a_52052_20860.t15 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X361 a_50583_13108.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X362 a_65534_25280# a_65088_25280# a_65438_25280# gnd sky130_fd_pr__nfet_01v8 ad=1.29323e+11p pd=1.01538e+06u as=5.94e+10p ps=690000u w=360000u l=150000u
X363 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X364 a_27962_11501# a_27762_11446.t13 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X365 Vso4b a_38070_8852.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X366 a_52052_20224# a_56272_15934.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X367 gnd gnd vinit.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X368 a_14266_8900.t0 a_25099_11445.t15 a_26016_10878.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X369 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X370 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X371 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X372 a_28994_5597# a_26036_4988.t15 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X373 Vso5b a_14910_6932.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X374 a_26589_11500# a_25099_11445.t16 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X375 a_55602_11692# a_51041_13108# a_52052_20860.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X376 gnd gnd vinit.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X377 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X378 a_26589_11500# a_25099_11445.t17 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X379 a_23919_5596# a_14188_14050.t18 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X380 a_24177_5596# a_14188_14050.t19 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X381 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X382 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X383 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X384 Fvco_By4_QPH_bar.t0 a_66167_26022# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X385 a_23160_10936.t5 a_14266_8900.t26 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X386 a_27962_11501# a_27762_11446.t14 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X387 a_77586_24654# a_77560_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X388 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X389 vinit.t12 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X390 a_64230_26048# RESET gnd gnd sky130_fd_pr__nfet_01v8 ad=6.405e+10p pd=725000u as=9.2007e+10p ps=682276u w=420000u l=150000u
X391 a_56602_11692# a_51636_13108# a_52052_20860.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X392 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X393 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X394 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X395 a_27962_11501# a_27762_11446.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X396 gnd gnd vbiasr.t14 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X397 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X398 a_28478_17218# a_26368_16652.t19 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X399 a_30384_802.t1 a_26036_4988.t16 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X400 z.t5 a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X401 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X402 a_4314_12044# a_4226_11996# a_4314_11948# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X403 a_26589_17217# a_23436_16644.t13 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X404 a_22629_17217# Fvco.t17 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X405 a_27962_11501# a_27762_11446.t16 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X406 gnd CLK_BY_2_BAR a_64911_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X407 a_65656_25522# a_65438_25280# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.27872e+11p pd=1.2608e+06u as=1.40201e+11p ps=1.03966e+06u w=640000u l=150000u
X408 a_28478_17218# a_26368_16652.t20 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X409 a_26073_5596# a_23414_5032.t15 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X410 zz CLK_BY_4_IPH_BAR.t3 a_34590_30714# vdd sky130_fd_pr__pfet_01v8 ad=6.012e+11p pd=4.62e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X411 a_22629_17217# Fvco.t18 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X412 a_23145_11500# a_14266_8900.t27 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X413 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X414 a_23160_10936.t4 a_14266_8900.t28 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X415 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X416 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X417 a_27962_17218# a_26368_16652.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X418 a_51041_13108# a_50511_16072.t8 a_50583_13108.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X419 a_66167_26022# RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X420 a_23160_10936.t3 a_14266_8900.t29 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X421 a_28220_11501# a_27762_11446.t17 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X422 a_28578_5014.t5 a_26036_4988.t17 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X423 a_57726_5786.t4 a_51532_4150.t4 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.72176e+11p ps=2.6849e+06u w=1.72e+06u l=4e+06u
X424 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X425 a_23160_10936.t2 a_14266_8900.t30 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X426 a_26847_17217# a_23436_16644.t14 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X427 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X428 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X429 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X430 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X431 a_63311_26048# a_62961_26048# a_63216_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.245e+10p pd=765000u as=6.51e+10p ps=730000u w=420000u l=150000u
X432 a_55602_11692# a_51041_13108# a_52052_20860.t13 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X433 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X434 a_65088_25280# a_64922_25280# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X435 a_23403_5596# a_14188_14050.t20 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X436 vdd a_54410_8156# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X437 a_23178_16644# Fvco.t19 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X438 CLK_IN a_23308_802.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X439 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X440 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X441 vinit.t34 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X442 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X443 a_50128_8156# a_54448_7822.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X444 a_65546_25646# a_64922_25280# a_65438_25280# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=7.245e+10p ps=765000u w=420000u l=150000u
X445 gnd a_17685_3840.t32 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X446 a_53308_2992# a_49874_4150.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.9575e+11p pd=1.64e+06u as=2.95737e+11p ps=2.19303e+06u w=1.35e+06u l=8e+06u
X447 gnd a_17685_3840.t33 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X448 a_28578_5014.t4 a_26036_4988.t18 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X449 vinit.t11 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X450 gnd Vso2b a_8736_14034# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X451 a_27962_5597# a_26036_4988.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X452 vdd a_4226_11996# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X453 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X454 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X455 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X456 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X457 gnd a_17685_3840.t34 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X458 Fvco.t0 a_26036_4988.t20 a_28578_5014.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X459 a_22629_5596# a_14188_14050.t21 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X460 a_26016_10878.t5 a_25099_11445.t18 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X461 a_25299_11500# a_25099_11445.t19 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X462 a_29510_5597# a_26036_4988.t21 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X463 a_23403_5596# a_14188_14050.t22 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X464 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X465 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X466 a_17685_3840.t4 vinit.t40 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=1e+06u
X467 a_23661_5596# a_14188_14050.t23 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X468 vinit.t10 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X469 vdd a_63876_26048# a_64051_26022# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X470 a_25299_11500# a_25099_11445.t20 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X471 a_23919_5596# a_14188_14050.t24 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X472 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X473 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X474 gnd a_17685_3840.t35 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X475 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X476 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X477 a_26073_11500# a_25099_11445.t21 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X478 vbiasr.t13 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X479 a_65077_26048# a_64911_26048# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.38484e+11p ps=999033u w=640000u l=150000u
X480 a_25299_17217# a_23436_16644.t15 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X481 Vso7b a_26690_784.t2 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X482 a_30384_802.t0 a_26036_4988.t22 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X483 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X484 a_26016_10878.t4 a_25099_11445.t22 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X485 a_25815_5596# a_23414_5032.t16 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X486 a_28736_5597# a_26036_4988.t23 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X487 a_26016_10878.t3 a_25099_11445.t23 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X488 a_29252_5597# a_26036_4988.t24 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X489 a_29510_5597# a_26036_4988.t25 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X490 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X491 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X492 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X493 a_66112_25280# a_64922_25280# a_66003_25280# gnd sky130_fd_pr__nfet_01v8 ad=6.17538e+10p pd=692308u as=7.11e+10p ps=755000u w=360000u l=150000u
X494 a_26016_10878.t2 a_25099_11445.t24 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X495 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X496 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X497 gnd a_17685_3840.t36 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X498 a_26073_11500# a_25099_11445.t25 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X499 vbiasr.t36 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X500 a_56602_11692# Fvco_By4_QPH_bar.t3 a_50320_14126# gnd sky130_fd_pr__nfet_01v8 ad=1.98421e+11p pd=1.49053e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X501 a_23156_5032.t6 a_14188_14050.t25 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X502 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X503 gnd a_17685_3840.t37 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X504 a_46856_21176.t1 a_51138_21494.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X505 gnd a_17685_3840.t38 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X506 a_26110_16652# a_23436_16644.t16 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X507 a_25557_17217# a_23436_16644.t17 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X508 a_26073_11500# a_25099_11445.t26 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X509 a_65645_26290# a_65427_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.27872e+11p pd=1.2608e+06u as=1.40201e+11p ps=1.03966e+06u w=640000u l=150000u
X510 a_26589_17217# a_23436_16644.t18 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X511 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X512 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X513 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X514 a_26073_11500# a_25099_11445.t27 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X515 a_26589_17217# a_23436_16644.t19 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X516 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X517 a_25815_5596# a_23414_5032.t17 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X518 vdd vdd vinit.t33 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X519 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X520 a_27962_17218# a_26368_16652.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X521 a_25557_5596# a_23414_5032.t18 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X522 a_42574_15624# vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=4e+06u
X523 gnd a_56334_20860.t2 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X524 a_26073_5596# a_23414_5032.t19 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X525 a_28478_5597# a_26036_4988.t26 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X526 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X527 gnd a_64051_26022# a_64615_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X528 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X529 a_29252_5597# a_26036_4988.t27 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X530 a_26073_17217# a_23436_16644.t20 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X531 a_24177_17217# Fvco.t20 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X532 a_27962_17218# a_26368_16652.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X533 a_77586_24654# CLK_BY_4_IPH_BAR.t0 gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X534 a_25778_4988.t5 a_23414_5032.t20 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X535 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X536 gnd a_17685_3840.t39 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X537 a_26331_11500# a_25099_11445.t28 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X538 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X539 gnd gnd vinit.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X540 vdd vinit.t41 a_17685_3840.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.16382e+11p pd=1.56099e+06u as=0p ps=0u w=1e+06u l=1e+06u
X541 a_28578_5014.t3 a_26036_4988.t28 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X542 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X543 a_65077_26048# a_64911_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X544 vbiasr.t12 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X545 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X546 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X547 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X548 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X549 vdd Vso3b a_4288_12110# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X550 a_77560_23350# a_77242_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X551 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X552 vdd CLK_BY_2_BAR a_64725_25280# vdd sky130_fd_pr__pfet_01v8_hvt ad=2.16382e+11p pd=1.56099e+06u as=1.35e+11p ps=1.27e+06u w=1e+06u l=150000u
X553 vdd Vso5b a_4288_11918# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X554 a_23178_16644# Fvco.t21 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X555 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X556 Vso3b a_32948_24994.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X557 a_25815_11500# a_25099_11445.t29 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X558 a_23403_5596# a_14188_14050.t26 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X559 a_23178_16644# Fvco.t22 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X560 a_25557_5596# a_23414_5032.t21 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X561 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X562 gnd gnd vinit.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X563 a_23504_23306# vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X564 a_25299_5596# a_23414_5032.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X565 a_51636_13108# a_50511_16072.t9 a_46856_19268.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=2e+06u
X566 a_26847_5596# a_23414_5032.t23 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X567 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X568 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X569 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X570 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X571 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X572 a_25815_11500# a_25099_11445.t30 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X573 vdd vdd vbiasr.t35 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X574 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X575 bb Fvco_By4_QPH.t4 a_47968_16078# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X576 a_28220_5597# a_26036_4988.t29 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X577 vdd Vso7b a_4226_11612# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X578 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X579 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X580 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X581 a_29510_11501# a_27762_11446.t18 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X582 a_25815_11500# a_25099_11445.t31 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X583 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X584 a_29510_5597# a_26036_4988.t30 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X585 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X586 a_25815_11500# a_25099_11445.t32 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X587 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X588 a_47968_16078# Fvco_By4_QPH_bar.t4 aa vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X589 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X590 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X591 a_25299_5596# a_23414_5032.t24 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X592 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X593 vdd vdd vbiasr.t34 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X594 Vso3b a_32948_24994.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X595 vdd Vso7b a_4288_11726# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X596 a_25815_17217# a_23436_16644.t21 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X597 a_25299_17217# a_23436_16644.t22 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X598 a_26589_5596# a_23414_5032.t25 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X599 a_23919_17217# Fvco.t23 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X600 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X601 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X602 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X603 a_25299_17217# a_23436_16644.t23 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X604 a_29510_11501# a_27762_11446.t19 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X605 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X606 a_25815_5596# a_23414_5032.t26 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X607 vinit.t32 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X608 a_63407_26048# a_62961_26048# a_63311_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.29323e+11p pd=1.01538e+06u as=5.94e+10p ps=690000u w=360000u l=150000u
X609 a_29510_11501# a_27762_11446.t20 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X610 CLK_IN a_23308_802.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X611 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X612 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X613 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X614 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X615 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X616 a_66101_26048# a_64911_26048# a_65992_26048# gnd sky130_fd_pr__nfet_01v8 ad=6.17538e+10p pd=692308u as=7.11e+10p ps=755000u w=360000u l=150000u
X617 a_25099_11445.t0 a_27762_11446.t21 a_28438_10874.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X618 a_28790_25040.t1 a_26368_16652.t24 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X619 a_22887_17217# Fvco.t24 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X620 a_29510_11501# a_27762_11446.t22 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X621 a_29252_5597# a_26036_4988.t31 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X622 a_65535_26414# RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=9.08803e+10p ps=655615u w=420000u l=150000u
X623 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X624 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X625 vinit.t7 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X626 a_26110_16652# a_23436_16644.t24 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X627 Vso5b a_14910_6932.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X628 a_23436_16644.t1 Fvco.t4 a_17685_3840.t15 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X629 vbiasot vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=4e+06u
X630 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X631 a_29510_17218# a_26368_16652.t25 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X632 Vso7b a_26690_784.t3 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X633 a_26110_16652# a_23436_16644.t25 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X634 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X635 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X636 a_23661_11500# a_14266_8900.t31 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X637 a_26073_17217# a_23436_16644.t26 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X638 a_25557_5596# a_23414_5032.t27 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X639 vdd Vso8b a_4288_11534# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X640 a_26331_5596# a_23414_5032.t28 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X641 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X642 gnd a_17685_3840.t40 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X643 a_26073_17217# a_23436_16644.t27 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X644 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X645 gnd a_17685_3840.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X646 a_50262_14152# Fvco_By4_QPH.t5 a_51041_13108# gnd sky130_fd_pr__nfet_01v8 ad=2.07143e+11p pd=1.67714e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X647 a_47968_16078# a_42550_16062# a_50511_16072.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X648 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X649 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X650 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X651 CLK_BY_2 a_64051_26022# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.8e+11p pd=2.56e+06u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X652 a_23145_11500# a_14266_8900.t32 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X653 a_49874_4150.t3 a_51532_4150.t5 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=3.59194e+11p ps=2.59124e+06u w=1.66e+06u l=4e+06u
X654 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X655 vdd CLK_IN a_4226_11420# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X656 vbiasr.t33 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X657 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X658 bb vbiasbuffer.t3 a_51826_16054.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=1e+06u
X659 a_28220_11501# a_27762_11446.t23 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X660 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X661 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.0669e+12p pd=2.27425e+07u as=3.0669e+12p ps=2.27425e+07u w=1.4e+07u l=1e+06u
X662 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X663 vinit.t31 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X664 a_28438_10874.t4 a_27762_11446.t24 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X665 a_43010_16058# Fvco_By4_QPH.t6 a_42574_15624# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X666 a_25299_5596# a_23414_5032.t29 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X667 Fvco_By4_QPH.t1 a_66731_26048# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X668 a_28994_11501# a_27762_11446.t25 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X669 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X670 a_23145_11500# a_14266_8900.t33 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X671 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X672 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X673 a_22629_17217# Fvco.t25 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X674 a_28994_11501# a_27762_11446.t26 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X675 a_23145_11500# a_14266_8900.t34 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X676 a_28220_11501# a_27762_11446.t27 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X677 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X678 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X679 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X680 a_23145_11500# a_14266_8900.t35 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X681 a_50511_16072.t4 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X682 vdd vdd vinit.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X683 a_66165_25646# a_65088_25280# a_66003_25280# vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=5.88e+10p ps=700000u w=420000u l=150000u
X684 a_28220_11501# a_27762_11446.t28 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X685 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X686 a_64051_26022# RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X687 a_65427_26048# a_65077_26048# a_65332_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=7.245e+10p pd=765000u as=6.51e+10p ps=730000u w=420000u l=150000u
X688 a_17685_3840.t2 vinit.t42 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=1e+06u
X689 a_23145_17217# Fvco.t4 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X690 a_28994_17218# a_26368_16652.t26 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X691 a_28220_11501# a_27762_11446.t29 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X692 a_42782_16060# vbiasot gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=4e+06u
X693 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X694 vdd a_51138_19904.t1 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X695 a_25815_17217# a_23436_16644.t28 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X696 a_23403_11500# a_14266_8900.t36 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X697 a_28220_17218# a_26368_16652.t27 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X698 a_25815_17217# a_23436_16644.t29 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X699 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X700 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X701 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X702 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X703 a_65992_26048# a_64911_26048# a_65645_26290# vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=8.61e+10p ps=790000u w=420000u l=150000u
X704 a_52052_20224# a_56334_19906# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X705 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X706 a_28994_17218# a_26368_16652.t28 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X707 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X708 a_24177_5596# a_14188_14050.t27 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X709 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X710 a_42550_16062# Fvco_By4_QPH.t7 a_42574_15624# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X711 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X712 a_23436_16644.t0 Fvco.t26 a_23178_16644# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X713 vbiasr.t32 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X714 a_77586_24654# a_77560_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X715 vdd vdd vinit.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X716 a_29510_17218# a_26368_16652.t29 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X717 a_22629_5596# a_14188_14050.t28 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X718 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X719 a_66003_25280# a_65088_25280# a_65656_25522# gnd sky130_fd_pr__nfet_01v8 ad=7.11e+10p pd=755000u as=7.1928e+10p ps=709200u w=360000u l=150000u
X720 Vso6b a_14832_12082.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X721 a_28736_11501# a_27762_11446.t30 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X722 gnd a_17685_3840.t42 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X723 a_4314_11660# a_4226_11612# a_4314_11564# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X724 a_29510_17218# a_26368_16652.t30 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X725 gnd gnd vbiasr.t11 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X726 gnd a_17685_3840.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X727 a_65343_25280# CLK_BY_4_IPH_BAR.t4 gnd gnd sky130_fd_pr__nfet_01v8 ad=7.10769e+10p pd=802308u as=9.2007e+10p ps=682276u w=420000u l=150000u
X728 a_28736_11501# a_27762_11446.t31 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X729 a_23919_5596# a_14188_14050.t29 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X730 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X731 a_28478_11501# a_27762_11446.t32 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X732 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X733 vdd vdd vinit.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X734 a_24177_5596# a_14188_14050.t30 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X735 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X736 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X737 a_23414_5032.t1 a_14188_14050.t31 a_17685_3840.t12 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X738 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X739 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X740 vdd vinit.t43 a_17685_3840.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=2.16382e+11p pd=1.56099e+06u as=0p ps=0u w=1e+06u l=1e+06u
X741 a_28736_17218# a_26368_16652.t31 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X742 gnd a_17685_3840.t44 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X743 a_28736_5597# a_26036_4988.t32 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X744 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X745 gnd a_17685_3840.t45 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X746 gnd a_17685_3840.t46 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X747 a_9628_32967# CLK_BY_4_IPH.t3 vctrl gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=3.012e+11p ps=2.62e+06u w=1e+06u l=150000u
X748 a_26331_11500# a_25099_11445.t33 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X749 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X750 a_23156_5032.t5 a_14188_14050.t32 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X751 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X752 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X753 a_28736_17218# a_26368_16652.t32 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X754 a_27962_5597# a_26036_4988.t33 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X755 a_77268_24654# CLK_BY_4_IPH.t0 gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X756 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X757 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X758 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X759 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X760 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X761 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X762 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X763 a_4314_11756# a_4288_11726# a_4314_11660# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X764 a_28478_5597# a_26036_4988.t34 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X765 a_23145_5596# a_14188_14050.t33 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X766 a_26331_11500# a_25099_11445.t34 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X767 a_23661_5596# a_14188_14050.t34 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X768 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X769 a_25778_4988.t4 a_23414_5032.t30 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X770 gnd gnd vbiasr.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X771 a_28994_17218# a_26368_16652.t33 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X772 a_26331_11500# a_25099_11445.t35 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X773 a_28578_5014.t2 a_26036_4988.t35 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X774 z.t4 a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X775 a_23145_17217# Fvco.t27 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X776 a_23308_802.t1 Fvco.t28 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X777 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X778 a_28994_17218# a_26368_16652.t34 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X779 a_26331_11500# a_25099_11445.t36 a_26073_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X780 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X781 a_23145_17217# Fvco.t29 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X782 a_42782_16060# Fvco_By4_QPH_bar.t5 a_43010_16058# vdd sky130_fd_pr__pfet_01v8 ad=3.72857e+11p pd=2.82e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X783 a_27962_5597# a_26036_4988.t36 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X784 a_28220_17218# a_26368_16652.t35 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X785 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X786 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X787 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X788 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X789 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X790 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X791 a_65343_25280# CLK_BY_4_IPH_BAR.t5 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=6.51e+10p pd=730000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X792 CLK_BY_4_IPH a_66178_25254# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X793 a_26331_17217# a_23436_16644.t30 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X794 a_23403_5596# a_14188_14050.t35 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X795 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X796 a_23178_16644# Fvco.t30 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X797 a_28220_17218# a_26368_16652.t36 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X798 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X799 a_22887_5596# a_14188_14050.t36 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X800 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X801 gnd a_17685_3840.t47 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X802 a_23661_5596# a_14188_14050.t37 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X803 a_26847_5596# a_23414_5032.t31 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X804 vdd Vso8b a_4226_11612# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X805 a_24177_5596# a_14188_14050.t38 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X806 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X807 a_65992_26048# a_65077_26048# a_65645_26290# gnd sky130_fd_pr__nfet_01v8 ad=7.11e+10p pd=755000u as=7.1928e+10p ps=709200u w=360000u l=150000u
X808 a_28220_5597# a_26036_4988.t37 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X809 a_77268_24654# a_77242_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X810 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X811 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X812 a_65332_26048# Fvco_By4_QPH.t8 gnd gnd sky130_fd_pr__nfet_01v8 ad=7.10769e+10p pd=802308u as=9.2007e+10p ps=682276u w=420000u l=150000u
X813 vbiasr.t31 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X814 a_46856_19268.t1 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X815 a_23414_5032.t0 a_14188_14050.t39 a_23156_5032.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X816 a_22629_5596# a_14188_14050.t40 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X817 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X818 a_26847_11500# a_25099_11445.t37 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X819 a_29510_5597# a_26036_4988.t38 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X820 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X821 vdd Vso6b a_4288_11726# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X822 a_26073_5596# a_23414_5032.t32 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X823 a_46856_21176.t0 a_51138_20858# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X824 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X825 a_26847_11500# a_25099_11445.t38 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X826 a_28994_5597# a_26036_4988.t39 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X827 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X828 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X829 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X830 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X831 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X832 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X833 a_26589_11500# a_25099_11445.t39 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X834 a_51826_16054.t0 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X835 a_26589_5596# a_23414_5032.t33 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X836 a_26036_4988.t1 a_23414_5032.t14 a_25778_4988.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X837 a_28736_17218# a_26368_16652.t37 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X838 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X839 gnd a_56334_20860.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X840 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X841 a_26847_17217# a_23436_16644.t31 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X842 a_28736_17218# a_26368_16652.t38 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X843 a_14266_8900.t1 a_25099_11445.t40 a_17685_3840.t14 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X844 a_23661_11500# a_14266_8900.t37 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X845 a_25815_5596# a_23414_5032.t34 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X846 a_51636_13108# Fvco_By4_QPH_bar.t6 a_51276_14152# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X847 a_28736_5597# a_26036_4988.t40 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X848 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X849 a_29252_5597# a_26036_4988.t41 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X850 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X851 vbiasr.t9 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X852 bb Fvco_By4_QPH.t9 a_47760_15642# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X853 a_26073_5596# a_23414_5032.t35 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X854 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X855 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X856 a_38070_8852.t0 a_25099_11445.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X857 vdd Vso2b a_4226_12188# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X858 a_23156_5032.t4 a_14188_14050.t41 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X859 a_26110_16652# a_23436_16644.t32 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X860 a_23661_11500# a_14266_8900.t38 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X861 a_27962_5597# a_26036_4988.t42 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X862 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X863 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X864 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X865 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X866 a_23661_11500# a_14266_8900.t39 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X867 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X868 a_28438_10874.t3 a_27762_11446.t33 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X869 a_26331_5596# a_23414_5032.t36 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X870 a_25557_5596# a_23414_5032.t37 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X871 a_55602_11692# Fvco_By4_QPH_bar.t7 a_50320_14126# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X872 gnd a_17685_3840.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X873 a_28478_5597# a_26036_4988.t43 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X874 a_23661_11500# a_14266_8900.t40 a_23403_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X875 vdd vdd vbiasr.t30 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X876 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X877 a_23661_5596# a_14188_14050.t42 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X878 vdd Vso3b a_4226_11996# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X879 a_26073_17217# a_23436_16644.t33 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X880 a_27762_11446.t1 a_26368_16652.t39 a_28622_16652# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.218e+11p ps=1.10264e+06u w=420000u l=1e+06u
X881 gnd a_17685_3840.t49 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X882 a_25778_4988.t3 a_23414_5032.t38 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X883 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X884 a_57726_5786.t1 a_57726_5786.t0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=6.57193e+11p ps=4.8734e+06u w=3e+06u l=1e+06u
X885 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X886 vdd a_65645_26290# a_65535_26414# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=1.134e+11p ps=1.1e+06u w=420000u l=150000u
X887 a_8752_10532# Vso7b a_4226_11612# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X888 a_23661_17217# Fvco.t4 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X889 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X890 aa Fvco_By4_QPH.t10 a_47968_16078# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X891 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X892 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X893 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X894 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X895 a_4314_12140# a_4288_12110# a_4314_12044# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X896 a_26331_17217# a_23436_16644.t34 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X897 a_28438_10874.t2 a_27762_11446.t34 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X898 vdd vdd vbiasr.t29 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X899 a_56602_11692# a_51636_13108# a_52052_20860.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X900 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X901 a_25557_11500# a_25099_11445.t42 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X902 a_62961_26048# a_62795_26048# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.38484e+11p ps=999033u w=640000u l=150000u
X903 gnd a_17685_3840.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X904 a_26331_17217# a_23436_16644.t35 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X905 a_28438_10874.t1 a_27762_11446.t35 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X906 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X907 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X908 zz CLK_BY_4_IPH_BAR.t6 a_9628_32967# gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X909 a_25557_11500# a_25099_11445.t43 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X910 Fvco.t1 a_26036_4988.t44 a_17685_3840.t16 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X911 a_25299_5596# a_23414_5032.t39 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X912 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X913 a_23403_11500# a_14266_8900.t41 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X914 a_28438_10874.t0 a_27762_11446.t36 a_29510_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X915 a_55602_11692# Fvco_By4_QPH_bar.t8 a_51334_14126# gnd sky130_fd_pr__nfet_01v8 ad=1.98421e+11p pd=1.49053e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X916 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X917 a_25299_11500# a_25099_11445.t44 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X918 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X919 vdd a_66178_25254# a_66742_25280# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X920 gnd gnd vbiasr.t8 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X921 a_26847_5596# a_23414_5032.t40 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X922 a_28622_16652# a_26368_16652.t40 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X923 a_25557_17217# a_23436_16644.t36 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X924 a_24177_11500# a_14266_8900.t42 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X925 a_28220_5597# a_26036_4988.t45 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X926 a_26690_784.t0 a_23414_5032.t41 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X927 a_29252_11501# a_27762_11446.t37 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X928 a_24177_11500# a_14266_8900.t43 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X929 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X930 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X931 a_23403_11500# a_14266_8900.t44 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X932 gnd gnd vbiasr.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X933 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X934 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X935 a_29252_11501# a_27762_11446.t38 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X936 a_55602_11692# a_51041_13108# a_52052_20860.t12 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X937 a_26073_5596# a_23414_5032.t42 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X938 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X939 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X940 a_23403_11500# a_14266_8900.t45 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X941 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X942 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X943 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X944 a_54966_3580# a_49874_4150.t9 a_53308_3580# gnd sky130_fd_pr__nfet_01v8 ad=7.0035e+11p pd=5.12e+06u as=7.0035e+11p ps=5.12e+06u w=4.83e+06u l=8e+06u
X945 vdd vdd vbiasr.t28 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X946 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X947 a_24177_17217# Fvco.t31 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X948 a_23403_11500# a_14266_8900.t46 a_23145_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X949 a_25815_17217# a_23436_16644.t37 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X950 a_47760_15642# Fvco_By4_QPH_bar.t9 bb vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.33143e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X951 a_26589_5596# a_23414_5032.t43 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X952 a_63216_26048# CLK_BY_2_BAR gnd gnd sky130_fd_pr__nfet_01v8 ad=7.10769e+10p pd=802308u as=9.2007e+10p ps=682276u w=420000u l=150000u
X953 a_26847_17217# a_23436_16644.t38 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X954 a_14188_14050.t1 a_14266_8900.t47 a_23160_10936.t7 gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X955 gnd a_4226_12188# a_4314_12140# gnd sky130_fd_pr__nfet_01v8 ad=7.09769e+11p pd=5.26327e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X956 vdd Vso5b a_4226_11804# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X957 a_29252_17218# a_26368_16652.t41 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X958 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X959 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X960 a_23403_17217# Fvco.t4 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X961 a_26847_17217# a_23436_16644.t39 a_26589_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X962 a_28478_11501# a_27762_11446.t39 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X963 a_51334_14126# Fvco_By4_QPH.t11 a_55602_11692# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X964 a_62961_26048# a_62795_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X965 vdd vdd vbiasr.t27 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X966 a_77560_23350# a_77242_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X967 vinit.t27 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X968 vbiasr.t26 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X969 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X970 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X971 vdd a_64051_26022# a_64615_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X972 gnd a_17685_3840.t51 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X973 vdd a_66178_25254# a_66165_25646# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X974 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X975 Vso2b a_28790_25040.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X976 a_65700_25280# a_65656_25522# a_65534_25280# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.50877e+11p ps=1.18462e+06u w=420000u l=150000u
X977 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X978 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X979 gnd gnd vinit.t6 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X980 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X981 a_29252_17218# a_26368_16652.t42 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X982 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X983 a_47760_15642# Fvco_By4_QPH_bar.t10 aa gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X984 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X985 a_22972_23306.t0 a_23504_23306# gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X986 a_28478_11501# a_27762_11446.t40 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X987 b a_77560_23350# gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X988 a_50262_14152# a_50320_14126# a_50511_16072.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X989 vdd CLK_IN a_62795_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X990 CLK_BY_4_IPH_BAR.t1 a_66742_25280# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X991 a_23919_11500# a_14266_8900.t48 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X992 a_28478_11501# a_27762_11446.t41 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X993 a_65535_26414# a_64911_26048# a_65427_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=7.245e+10p ps=765000u w=420000u l=150000u
X994 vdd a_54468_7504.t0 gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X995 a_23919_11500# a_14266_8900.t49 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X996 a_28478_11501# a_27762_11446.t42 a_28220_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X997 a_26331_5596# a_23414_5032.t44 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X998 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X999 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1000 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1001 a_23661_17217# Fvco.t32 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1002 vbiasr.t6 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1003 a_22887_11500# a_14266_8900.t50 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1004 a_47968_16078# Fvco_By4_QPH_bar.t11 bb gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1005 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1006 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1007 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1008 Vso1b a_24410_25128.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1009 a_28478_17218# a_26368_16652.t43 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1010 a_23661_17217# Fvco.t33 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1011 a_23919_17217# Fvco.t34 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1012 a_22887_11500# a_14266_8900.t51 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1013 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1014 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1015 a_42550_16062# Fvco_By4_QPH.t12 a_42782_16060# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=3.72857e+11p ps=2.82e+06u w=2e+06u l=150000u
X1016 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1017 vbiasr.t25 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1018 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1019 a_22887_17217# Fvco.t4 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1020 Vso4b a_38070_8852.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1021 a_52052_20860.t2 a_51636_13108# a_56602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X1022 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1023 CLK_BY_2 a_64051_26022# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.69e+11p pd=1.82e+06u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X1024 a_28622_16652# a_26368_16652.t44 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1025 a_23145_5596# a_14188_14050.t43 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1026 gnd RESET a_65700_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=4.41e+10p ps=630000u w=420000u l=150000u
X1027 gnd a_66178_25254# a_66112_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=7.20462e+10p ps=807692u w=420000u l=150000u
X1028 a_25557_17217# a_23436_16644.t40 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1029 a_51532_4150.t3 a_49932_4124.t3 a_49874_4150.t2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.28e+06u l=8e+06u
X1030 a_64725_25280# CLK_BY_2_BAR gnd gnd sky130_fd_pr__nfet_01v8 ad=8.775e+10p pd=920000u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X1031 vdd a_4288_11534# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1032 a_28622_16652# a_26368_16652.t45 a_29510_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1033 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1034 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1035 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1036 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1037 CLK_BY_4_IPH.t1 a_66178_25254# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X1038 a_17685_3840.t8 vctrl a_22972_23306.t3 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1039 a_25557_17217# a_23436_16644.t41 a_25299_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1040 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1041 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1042 vdd vdd vinit.t26 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1043 vinit.t5 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1044 gnd CLK_IN a_62795_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1045 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1046 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1047 a_23145_17217# Fvco.t35 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1048 a_24177_17217# Fvco.t36 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1049 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1050 gnd a_17685_3840.t52 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1051 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1052 a_9628_32967# CLK_BY_4_IPH.t4 zz vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=6.012e+11p ps=4.62e+06u w=2e+06u l=150000u
X1053 a_24177_17217# Fvco.t37 a_23919_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1054 vbiasr.t5 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1055 gnd a_17685_3840.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1056 vinit.t4 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1057 a_29252_17218# a_26368_16652.t46 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1058 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1059 a_65645_26290# a_65427_26048# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.722e+11p pd=1.58e+06u as=1.81761e+11p ps=1.31123e+06u w=840000u l=150000u
X1060 a_23403_17217# Fvco.t38 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1061 a_22887_5596# a_14188_14050.t44 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1062 a_52052_20860.t11 a_51041_13108# a_55602_11692# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=7.93684e+11p ps=5.96211e+06u w=4e+06u l=1e+06u
X1063 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1064 a_29252_17218# a_26368_16652.t47 a_28994_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1065 a_23403_17217# Fvco.t39 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1066 a_26589_11500# a_25099_11445.t45 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1067 a_22629_11500# a_14266_8900.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1068 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1069 a_24177_5596# a_14188_14050.t45 a_23919_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1070 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1071 a_34590_30714# CLK_BY_4_IPH.t5 zz gnd sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.33e+06u as=1.65e+11p ps=1.33e+06u w=1e+06u l=150000u
X1072 a_22629_11500# a_14266_8900.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1073 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1074 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1075 a_50511_16072.t6 a_42550_16062# a_47968_16078# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1076 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1077 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1078 vdd a_51138_20858# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1079 gnd a_17685_3840.t54 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1080 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1081 a_22629_17217# Fvco.t4 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1082 Fvco_By4_QPH.t0 a_66731_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.42392e+11p ps=1.0559e+06u w=650000u l=150000u
X1083 Vso6b a_14832_12082.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1084 vdd Vso4b a_4226_11996# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1085 a_26589_11500# a_25099_11445.t46 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1086 a_28994_5597# a_26036_4988.t46 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1087 a_56602_11692# a_51636_13108# a_52052_20860.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1088 a_50511_16072.t2 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1089 a_51276_14152# Fvco_By4_QPH.t13 a_51041_13108# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1090 a_26589_11500# a_25099_11445.t47 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1091 vdd vdd vinit.t25 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1092 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1093 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1094 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1095 a_26589_11500# a_25099_11445.t48 a_26331_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1096 vdd vdd vbiasr.t24 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1097 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1098 a_77586_24654# a_77560_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1099 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1100 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1101 a_28478_17218# a_26368_16652.t48 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1102 vdd Vso1b a_4226_12188# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1103 a_26589_17217# a_23436_16644.t42 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1104 a_23919_17217# Fvco.t40 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1105 a_28478_17218# a_26368_16652.t49 a_28220_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1106 a_28994_11501# a_27762_11446.t43 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1107 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.416e+07u w=2.4e+07u
X1108 a_56602_11692# Fvco_By4_QPH_bar.t12 a_51334_14126# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1109 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1110 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1111 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1112 vinit.t24 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1113 a_63419_26414# a_62795_26048# a_63311_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=7.245e+10p ps=765000u w=420000u l=150000u
X1114 a_23919_17217# Fvco.t41 a_23661_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1115 a_43010_16058# Fvco_By4_QPH.t14 a_42782_16060# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1116 a_55602_11692# a_51041_13108# a_52052_20860.t10 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1117 a_24410_25128.t0 a_23436_16644.t43 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1118 a_63876_26048# a_62795_26048# a_63529_26290# vdd sky130_fd_pr__pfet_01v8_hvt ad=5.88e+10p pd=700000u as=8.61e+10p ps=790000u w=420000u l=150000u
X1119 a_22887_17217# Fvco.t42 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1120 a_27962_5597# a_26036_4988.t47 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1121 a_53292_4814# a_49874_4150.t10 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.856e+11p pd=1.57e+06u as=2.80402e+11p ps=2.07932e+06u w=1.28e+06u l=8e+06u
X1122 gnd a_66167_26022# a_66101_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=7.20462e+10p ps=807692u w=420000u l=150000u
X1123 gnd RESET a_65689_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=4.41e+10p ps=630000u w=420000u l=150000u
X1124 a_22887_17217# Fvco.t43 a_22629_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1125 gnd a_17685_3840.t55 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1126 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1127 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1128 a_22629_5596# a_14188_14050.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1129 gnd a_17685_3840.t56 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1130 a_23145_5596# a_14188_14050.t47 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1131 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1132 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1133 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1134 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1135 a_63529_26290# a_63311_26048# gnd gnd sky130_fd_pr__nfet_01v8 ad=1.27872e+11p pd=1.2608e+06u as=1.40201e+11p ps=1.03966e+06u w=640000u l=150000u
X1136 a_23661_5596# a_14188_14050.t48 a_23403_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1137 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=3.0669e+12p pd=2.27425e+07u as=3.0669e+12p ps=2.27425e+07u w=1.4e+07u l=1e+06u
X1138 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=2.19064e+11p pd=1.62447e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1139 a_28790_25040.t0 a_26368_16652.t50 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1140 a_25299_11500# a_25099_11445.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1141 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1142 Vso8b a_30384_802.t2 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.218e+11p pd=1.42e+06u as=9.2007e+10p ps=682276u w=420000u l=150000u
X1143 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1144 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1145 vdd Vso2b a_4288_12110# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1146 a_46856_19268.t2 gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1147 vdd Vso4b a_4288_11918# vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1148 a_56602_11692# a_51636_13108# a_52052_20860.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1149 gnd a_17685_3840.t57 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1150 a_42782_16060# bb a_44752_16348.t4 vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1151 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1152 a_64051_26022# a_63876_26048# a_64230_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=6.405e+10p ps=725000u w=420000u l=150000u
X1153 a_8748_11114# Vso6b a_4288_11726# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1154 a_26331_17217# a_23436_16644.t44 a_26073_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1155 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1156 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1157 a_28736_5597# a_26036_4988.t48 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1158 a_22629_5596# a_14188_14050.t49 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1159 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1160 a_25299_11500# a_25099_11445.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1161 a_22887_5596# a_14188_14050.t50 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1162 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1163 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1164 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1165 a_25299_11500# a_25099_11445.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1166 a_23919_5596# a_14188_14050.t51 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1167 vinit.t23 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1168 a_28736_11501# a_27762_11446.t44 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1169 vbiasot a_51532_4150.t6 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.566e+11p pd=1.66e+06u as=1.16846e+11p ps=842934u w=540000u l=8e+06u
X1170 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1171 a_27962_11501# a_27762_11446.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1172 a_25299_11500# a_25099_11445.t52 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1173 a_23156_5032.t3 a_14188_14050.t52 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1174 vbiasbuffer.t2 vbiasbuffer.t1 a_54468_7504.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1175 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1176 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1177 a_14188_14050.t0 a_14266_8900.t54 a_17685_3840.t11 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1178 a_27962_11501# a_27762_11446.t46 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1179 a_55602_11692# a_51041_13108# a_52052_20860.t9 gnd sky130_fd_pr__nfet_01v8_lvt ad=7.93684e+11p pd=5.96211e+06u as=0p ps=0u w=4e+06u l=1e+06u
X1180 a_51334_14126# Fvco_By4_QPH.t15 a_56602_11692# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=1.98421e+11p ps=1.49053e+06u w=1e+06u l=150000u
X1181 a_25299_17217# a_23436_16644.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1182 a_22629_17217# Fvco.t44 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1183 gnd a_17685_3840.t58 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1184 a_42574_15624# aa a_44752_16348.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=9.32143e+11p pd=7.05e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1185 a_26073_5596# a_23414_5032.t45 a_25815_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1186 a_28736_5597# a_26036_4988.t49 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1187 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1188 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1189 a_24410_25128.t1 a_23436_16644.t46 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X1190 vdd a_4288_11726# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1191 a_14832_12082.t0 a_14188_14050.t53 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1192 a_22629_17217# Fvco.t45 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1193 a_28478_5597# a_26036_4988.t50 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1194 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1195 a_50128_8156# a_54410_8156# gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1196 a_28994_5597# a_26036_4988.t51 a_28736_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1197 a_23160_10936.t1 a_14266_8900.t55 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1198 a_42574_15624# Fvco_By4_QPH_bar.t13 a_43010_16058# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1199 a_17685_3840.t0 vinit.t44 vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=1e+06u
X1200 a_27962_17218# a_26368_16652.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1201 a_25778_4988.t2 a_23414_5032.t46 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1202 a_54966_2992# a_49874_4150.t11 a_53308_2992# gnd sky130_fd_pr__nfet_01v8 ad=1.9575e+11p pd=1.64e+06u as=1.9575e+11p ps=1.64e+06u w=1.35e+06u l=8e+06u
X1203 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1204 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1205 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1206 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1207 a_25099_11445.t1 a_27762_11446.t47 a_17685_3840.t13 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1208 a_23160_10936.t0 a_14266_8900.t56 a_24177_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1209 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1210 a_22972_23306.t2 vctrl a_17685_3840.t7 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1211 a_23156_5032.t2 a_14188_14050.t54 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1212 vctrl CLK_BY_4_IPH_BAR.t7 a_9628_32967# vdd sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.33e+06u as=3.3e+11p ps=2.33e+06u w=2e+06u l=150000u
X1213 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1214 a_17685_3840.t9 vctrl a_22972_23306.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=2e+06u
X1215 a_26589_17217# a_23436_16644.t47 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1216 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1217 a_8740_12844# Vso3b a_4226_11996# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1218 a_4314_11468# a_4226_11420# vout gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=1.0044e+12p ps=7.1e+06u w=3.24e+06u l=150000u
X1219 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1220 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1221 a_66154_26414# a_65077_26048# a_65992_26048# vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=5.88e+10p ps=700000u w=420000u l=150000u
X1222 a_27762_11446.t0 a_26368_16652.t52 a_17685_3840.t10 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1223 a_26589_17217# a_23436_16644.t48 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1224 a_38070_8852.t1 a_25099_11445.t53 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.1901e+11p ps=858544u w=550000u l=8e+06u
X1225 a a_77242_23350# gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X1226 a_23178_16644# Fvco.t46 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1227 a_27962_17218# a_26368_16652.t53 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1228 a_28478_5597# a_26036_4988.t52 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1229 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1230 a_22972_23306.t4 vdd gnd sky130_fd_pr__res_xhigh_po_0p35 l=500000u
X1231 a_51041_13108# Fvco_By4_QPH_bar.t14 a_50262_14152# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1232 a_25778_4988.t1 a_23414_5032.t47 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1233 a_26847_5596# a_23414_5032.t48 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1234 a_32948_24994.t0 a_27762_11446.t48 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=150000u
X1235 vbiasr.t23 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1236 a_28578_5014.t1 a_26036_4988.t53 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1237 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1238 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1239 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1240 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1241 a_63419_26414# RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.134e+11p pd=1.1e+06u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1242 a_28220_5597# a_26036_4988.t54 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1243 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1244 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1245 a_77268_24654# a_77242_23350# sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1246 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1247 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1248 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1249 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1250 a_22629_5596# a_14188_14050.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1251 a_55602_11692# vbiasob.t4 a_51138_21494.t0 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=2e+06u
X1252 a_23403_5596# a_14188_14050.t56 a_23145_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1253 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1254 vdd vdd vinit.t22 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1255 vdd a_4226_11612# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1256 a_23661_17217# Fvco.t47 a_23403_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1257 a_51041_13108# Fvco_By4_QPH_bar.t15 a_51276_14152# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.07143e+11p ps=1.67714e+06u w=1e+06u l=150000u
X1258 a_26847_5596# a_23414_5032.t49 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1259 a_26589_5596# a_23414_5032.t50 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1260 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1261 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1262 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1263 a_28220_5597# a_26036_4988.t55 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1264 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1265 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1266 vdd a_64051_26022# a_64038_26414# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X1267 a_4314_11852# a_4226_11804# a_4314_11756# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X1268 a_26016_10878.t1 a_25099_11445.t54 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1269 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1270 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1271 gnd a_66178_25254# a_66742_25280# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1272 a_26016_10878.t0 a_25099_11445.t55 a_26847_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1273 a_28736_5597# a_26036_4988.t56 a_28478_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1274 a_29510_5597# a_26036_4988.t57 a_29252_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1275 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1276 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1277 aa vbiasbuffer.t4 a_50032_16080.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.09667e+07u as=0p ps=0u w=5e+06u l=1e+06u
X1278 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1279 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1280 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1281 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1282 a_26847_11500# a_25099_11445.t56 a_26589_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1283 a_51636_13108# Fvco_By4_QPH_bar.t16 a_50262_14152# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.07143e+11p ps=1.67714e+06u w=1e+06u l=150000u
X1284 gnd gnd vinit.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1285 vdd a_66003_25280# a_66178_25254# vdd sky130_fd_pr__pfet_01v8_hvt ad=9.08803e+10p pd=655615u as=5.67e+10p ps=690000u w=420000u l=150000u
X1286 a_8748_11692# Vso5b a_4226_11804# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1287 a_26073_11500# a_25099_11445.t57 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1288 vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1289 a_50262_14152# Fvco_By4_QPH.t16 a_51636_13108# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=150000u
X1290 a_23156_5032.t1 a_14188_14050.t57 a_24177_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1291 CLK_BY_2_BAR a_64615_26048# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=2.6e+11p pd=2.52e+06u as=2.16382e+11p ps=1.56099e+06u w=1e+06u l=150000u
X1292 a_8744_9386# CLK_IN a_4226_11420# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1293 gnd a_17685_3840.t59 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1294 a_26589_5596# a_23414_5032.t51 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1295 a_26110_16652# a_23436_16644.t49 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1296 a_25299_17217# a_23436_16644.t50 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1297 a_26073_11500# a_25099_11445.t58 a_25815_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1298 a_65427_26048# a_64911_26048# a_65332_26048# gnd sky130_fd_pr__nfet_01v8 ad=5.94e+10p pd=690000u as=6.09231e+10p ps=687692u w=360000u l=150000u
X1299 vdd a_64725_25280# a_64922_25280# vdd sky130_fd_pr__pfet_01v8_hvt ad=1.38484e+11p pd=999033u as=1.664e+11p ps=1.8e+06u w=640000u l=150000u
X1300 a_25299_17217# a_23436_16644.t51 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1301 gnd a_17685_3840.t60 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1302 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1303 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1304 gnd gnd vbiasr.t4 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1305 a_44752_16348.t3 bb a_42782_16060# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1306 a_25815_5596# a_23414_5032.t52 a_25557_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1307 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1308 a_27962_17218# a_26368_16652.t54 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1309 a_26331_5596# a_23414_5032.t53 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1310 gnd a_17685_3840.t61 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1311 a_28478_5597# a_26036_4988.t58 a_28220_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1312 a_66178_25254# a_66003_25280# a_66357_25280# gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=6.405e+10p ps=725000u w=420000u l=150000u
X1313 gnd Vso8b a_8752_10532# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1314 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1315 a_29252_5597# a_26036_4988.t59 a_28994_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1316 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1317 a_26073_17217# a_23436_16644.t52 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1318 a_27962_17218# a_26368_16652.t55 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1319 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X1320 a_25778_4988.t0 a_23414_5032.t54 a_26847_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1321 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1322 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1323 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1324 a_47760_15642# a_43010_16058# z.t1 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.45e+12p pd=1.08286e+07u as=0p ps=0u w=5e+06u l=1e+06u
X1325 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1326 a_63529_26290# a_63311_26048# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.722e+11p pd=1.58e+06u as=1.81761e+11p ps=1.31123e+06u w=840000u l=150000u
X1327 a_23403_17217# Fvco.t48 a_23145_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1328 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1329 a_4314_11948# a_4288_11918# a_4314_11852# gnd sky130_fd_pr__nfet_01v8 ad=5.346e+11p pd=3.57e+06u as=5.346e+11p ps=3.57e+06u w=3.24e+06u l=150000u
X1330 gnd a_17685_3840.t62 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1331 a_23178_16644# Fvco.t49 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1332 a_51532_4150.t2 a_49874_4150.t12 a_54966_3580# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.0035e+11p ps=5.12e+06u w=4.83e+06u l=8e+06u
X1333 gnd CLK_BY_2_BAR a_64725_25280# gnd sky130_fd_pr__nfet_01v8 ad=1.42392e+11p pd=1.0559e+06u as=8.775e+10p ps=920000u w=650000u l=150000u
X1334 a_23178_16644# Fvco.t50 a_24177_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1335 a_25557_5596# a_23414_5032.t55 a_25299_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1336 a_44752_16348.t0 aa a_42574_15624# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=9.32143e+11p ps=7.05e+06u w=5e+06u l=1e+06u
X1337 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1338 a_26331_5596# a_23414_5032.t56 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1339 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1340 gnd Vso6b a_8748_11692# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1341 a_28994_11501# a_27762_11446.t49 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1342 a_26847_5596# a_23414_5032.t57 a_26589_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1343 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1344 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1345 a_65332_26048# Fvco_By4_QPH.t17 vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=6.51e+10p pd=730000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1346 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1347 vbiasr.t22 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1348 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1349 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1350 a_25815_11500# a_25099_11445.t59 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1351 a_28220_5597# a_26036_4988.t60 a_27962_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1352 a_25815_11500# a_25099_11445.t60 a_25557_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1353 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1354 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1355 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1356 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1357 a_8748_9956# Vso8b a_4288_11534# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1358 gnd a_17685_3840.t63 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1359 a_25557_11500# a_25099_11445.t61 a_25299_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1360 vinit.t2 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1361 a_28994_11501# a_27762_11446.t50 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1362 a_25299_5596# a_23414_5032.t58 gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=2.19064e+11p ps=1.62447e+06u w=1e+06u l=1e+06u
X1363 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1364 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1365 a_66178_25254# RESET vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=5.67e+10p pd=690000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1366 a_28994_11501# a_27762_11446.t51 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1367 gnd gnd vbiasr.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1368 vdd a_4288_12110# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1369 a_25815_17217# a_23436_16644.t53 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1370 a_26589_5596# a_23414_5032.t59 a_26331_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1371 vinit.t21 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1372 a_28994_11501# a_27762_11446.t52 a_28736_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1373 Vso8b a_30384_802.t3 vdd vdd sky130_fd_pr__pfet_01v8 ad=4.872e+11p pd=3.94e+06u as=3.63521e+11p ps=2.62246e+06u w=1.68e+06u l=150000u
X1374 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1375 gnd a_66167_26022# a_66731_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=1.092e+11p ps=1.36e+06u w=420000u l=150000u
X1376 a_29510_11501# a_27762_11446.t53 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1377 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.413e+07u w=2.4e+07u
X1378 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1379 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1380 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1381 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1382 a_24177_11500# a_14266_8900.t57 a_23919_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1383 vbiasr.t2 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1384 z.t0 a_43010_16058# a_47760_15642# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.45e+12p ps=1.08286e+07u w=5e+06u l=1e+06u
X1385 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1386 a_29510_11501# a_27762_11446.t54 a_29252_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1387 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1388 a_28994_17218# a_26368_16652.t56 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1389 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1390 gnd a_17685_3840.t64 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.53345e+12p pd=1.13713e+07u as=1.53345e+12p ps=1.13713e+07u w=7e+06u l=8e+06u
X1391 a_29252_11501# a_27762_11446.t55 a_28994_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1392 gnd gnd gnd sky130_fd_pr__res_xhigh_po w=350000u l=2.363e+07u
X1393 a_42782_16060# Fvco_By4_QPH_bar.t17 a_42550_16062# gnd sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1394 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1395 gnd a_64051_26022# a_63985_26048# gnd sky130_fd_pr__nfet_01v8 ad=9.2007e+10p pd=682276u as=7.20462e+10p ps=807692u w=420000u l=150000u
X1396 a_26110_16652# a_23436_16644.t54 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1397 a_50320_14126# Fvco_By4_QPH.t18 a_56602_11692# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.38667e+06u w=2e+06u l=150000u
X1398 a_29510_17218# a_26368_16652.t57 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1399 a_63985_26048# a_62795_26048# a_63876_26048# gnd sky130_fd_pr__nfet_01v8 ad=6.17538e+10p pd=692308u as=7.11e+10p ps=755000u w=360000u l=150000u
X1400 a_26110_16652# a_23436_16644.t55 a_26847_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.62534e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1401 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1402 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1403 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1404 a_28736_11501# a_27762_11446.t56 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1405 a_50262_14152# a_50320_14126# a_50511_16072.t1 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X1406 a_66167_26022# a_65992_26048# a_66346_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.092e+11p pd=1.36e+06u as=6.405e+10p ps=725000u w=420000u l=150000u
X1407 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1408 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1409 a_26073_17217# a_23436_16644.t56 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1410 a_51276_14152# a_51334_14126# z.t3 gnd sky130_fd_pr__nfet_01v8_lvt ad=4.14286e+11p pd=3.35429e+06u as=0p ps=0u w=2e+06u l=1e+06u
X1411 gnd gnd sky130_fd_pr__cap_mim_m3_1 l=2.41e+07u w=2.4e+07u
X1412 a_26331_5596# a_23414_5032.t60 a_26073_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1413 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1414 a_26073_17217# a_23436_16644.t57 a_25815_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1415 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1416 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1417 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1418 vinit.t1 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1419 vdd a_4226_11804# vout vdd sky130_fd_pr__pfet_01v8 ad=3.63521e+11p pd=2.62246e+06u as=4.872e+11p ps=3.94e+06u w=1.68e+06u l=150000u
X1420 a_29510_17218# a_26368_16652.t58 a_29252_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1421 a_28736_11501# a_27762_11446.t57 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1422 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1423 a_65088_25280# a_64922_25280# vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=1.664e+11p pd=1.8e+06u as=1.38484e+11p ps=999033u w=640000u l=150000u
X1424 a_28736_11501# a_27762_11446.t58 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1425 a_23919_5596# a_14188_14050.t58 a_23661_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1426 a_50511_16072.t0 a_50320_14126# a_50262_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1427 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1428 a_28736_11501# a_27762_11446.t59 a_28478_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1429 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1430 gnd gnd vinit.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1431 a_23919_11500# a_14266_8900.t58 a_23661_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1432 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1433 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1434 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1435 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1436 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1437 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1438 a_8736_14034# Vso1b a_4226_12188# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1439 vbiasr.t1 gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.09532e+12p ps=8.12233e+06u w=5e+06u l=1e+06u
X1440 a_65689_26048# a_65645_26290# a_65523_26048# gnd sky130_fd_pr__nfet_01v8 ad=4.41e+10p pd=630000u as=1.50877e+11p ps=1.18462e+06u w=420000u l=150000u
X1441 a_28736_17218# a_26368_16652.t59 a_28478_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1442 a_23145_11500# a_14266_8900.t59 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1443 a_23145_5596# a_14188_14050.t59 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1444 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1445 a_63876_26048# a_62961_26048# a_63529_26290# gnd sky130_fd_pr__nfet_01v8 ad=7.11e+10p pd=755000u as=7.1928e+10p ps=709200u w=360000u l=150000u
X1446 a_23145_11500# a_14266_8900.t60 a_22887_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1447 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1448 gnd gnd gnd sky130_fd_pr__res_xhigh_po_0p35 l=1.925e+07u
X1449 a_65523_26048# a_65077_26048# a_65427_26048# gnd sky130_fd_pr__nfet_01v8 ad=1.29323e+11p pd=1.01538e+06u as=5.94e+10p ps=690000u w=360000u l=150000u
X1450 gnd CLK_IN a_8748_9956# gnd sky130_fd_pr__nfet_01v8 ad=1.62108e+11p pd=1.2021e+06u as=1.221e+11p ps=1.07e+06u w=740000u l=150000u
X1451 a_28220_11501# a_27762_11446.t60 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1452 gnd gnd vbiasr.t0 gnd sky130_fd_pr__nfet_01v8_lvt ad=1.09532e+12p pd=8.12233e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1453 a_22887_11500# a_14266_8900.t61 a_22629_11500# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1454 a_28220_11501# a_27762_11446.t61 a_27962_11501# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1455 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1456 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1457 a_23145_17217# Fvco.t4 a_22887_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1458 a_63216_26048# CLK_BY_2_BAR vdd vdd sky130_fd_pr__pfet_01v8_hvt ad=6.51e+10p pd=730000u as=9.08803e+10p ps=655615u w=420000u l=150000u
X1459 a_25815_17217# a_23436_16644.t58 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1460 z.t2 a_51334_14126# a_51276_14152# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.14286e+11p ps=3.35429e+06u w=2e+06u l=1e+06u
X1461 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1462 a_28220_17218# a_26368_16652.t60 a_27962_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1463 a_26589_17217# a_23436_16644.t59 a_26331_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1464 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1465 a_26368_16652.t0 a_23436_16644.t60 a_17685_3840.t5 vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=4e+06u
X1466 a_25815_17217# a_23436_16644.t61 a_25557_17217# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1467 a_23145_5596# a_14188_14050.t60 a_22887_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1468 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1469 a_8744_13422# Vso2b a_4288_12110# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1470 a_22887_5596# a_14188_14050.t61 a_22629_5596# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1471 vdd vdd vbiasr.t21 vdd sky130_fd_pr__pfet_01v8_lvt ad=1.08191e+12p pd=7.80494e+06u as=0p ps=0u w=5e+06u l=1e+06u
X1472 aa Fvco_By4_QPH.t19 a_47760_15642# vdd sky130_fd_pr__pfet_01v8 ad=5.8e+11p pd=4.38667e+06u as=5.8e+11p ps=4.33143e+06u w=2e+06u l=150000u
X1473 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1474 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1475 vdd a_9628_32967# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1476 vinit.t20 vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.08191e+12p ps=7.80494e+06u w=5e+06u l=1e+06u
X1477 a_8748_12270# Vso4b a_4288_11918# gnd sky130_fd_pr__nfet_01v8 ad=1.221e+11p pd=1.07e+06u as=2.294e+11p ps=2.1e+06u w=740000u l=150000u
X1478 vdd a_34590_30714# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.51467e+12p pd=1.09269e+07u as=1.51467e+12p ps=1.09269e+07u w=7e+06u l=8e+06u
X1479 a_28994_17218# a_26368_16652.t61 a_28736_17218# gnd sky130_fd_pr__nfet_01v8_lvt ad=1.45e+11p pd=1.29e+06u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
X1480 a_28578_5014.t0 a_26036_4988.t61 a_29510_5597# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.45e+11p ps=1.29e+06u w=1e+06u l=1e+06u
C0 a_51636_13108# a_56602_11692# 2.40fF
C1 a_51334_14126# a_55602_11692# 2.35fF
C2 a_51276_14152# a_51041_13108# 2.50fF
C3 a_77586_24654# a_77268_24654# 10.04fF
C4 Vso2b Vso1b 3.79fF
C5 Fvco_By4_QPH_bar bb 2.30fF
C6 a_42550_16062# a_43010_16058# 4.58fF
C7 vdd a_4226_11996# 2.88fF
C8 vdd a_4288_11726# 2.30fF
C9 a_56602_11692# a_50320_14126# 2.53fF
C10 vdd Vso7b 2.92fF
C11 a_77560_23350# a_77586_24654# 155.27fF
C12 a_42550_16062# a_42782_16060# 2.13fF
C13 a_51334_14126# z 3.18fF
C14 a_42574_15624# a_43010_16058# 2.25fF
C15 a_9628_32967# vdd 505.89fF
C16 vbiasob vdd 2.62fF
C17 vinit vdd 36.67fF
C18 a_42550_16062# vdd 2.55fF
C19 a_55602_11692# a_50320_14126# 2.15fF
C20 bb a_47760_15642# 4.36fF
C21 vdd CLK_BY_4_IPH 5.66fF
C22 a_77560_23350# a_77268_24654# 14.35fF
C23 a_42574_15624# a_42782_16060# 2.88fF
C24 a_4226_12188# vout 2.67fF
C25 Vso2b vdd 3.24fF
C26 a_47968_16078# aa 3.02fF
C27 a_4226_11804# vdd 2.43fF
C28 vdd Vso3b 3.96fF
C29 a_51334_14126# a_50320_14126# 2.95fF
C30 a_77242_23350# a_77586_24654# 3.69fF
C31 vout vdd 7.94fF
C32 a_50262_14152# a_51636_13108# 2.25fF
C33 a_51276_14152# a_51636_13108# 2.56fF
C34 a_77242_23350# a_77268_24654# 117.99fF
C35 vdd a_4288_12110# 2.60fF
C36 Fvco_By4_QPH_bar Fvco_By4_QPH 16.00fF
C37 CLK_IN Vso4b 26.23fF
C38 vdd Vso5b 5.20fF
C39 RESET Fvco_By4_QPH 2.21fF
C40 vdd a_4226_11420# 2.26fF
C41 Vso8b Vso7b 12.19fF
C42 vdd Vso6b 3.09fF
C43 vctrl Vso1b 3.89fF
C44 a_42550_16062# a_42574_15624# 2.35fF
C45 Vso1b vdd 3.70fF
C46 a_77560_23350# a_77242_23350# 62.20fF
C47 a_55602_11692# a_56602_11692# 2.04fF
C48 a_47760_15642# a_47968_16078# 3.20fF
C49 vdd a_4288_11918# 2.56fF
C50 Vso4b vdd 3.85fF
C51 a_42782_16060# a_43010_16058# 2.44fF
C52 a_51041_13108# a_51636_13108# 4.40fF
C53 a_34590_30714# vdd 504.98fF
C54 bb a_47968_16078# 2.43fF
C55 a_4226_11612# vdd 2.37fF
C56 a_47760_15642# aa 2.29fF
C57 vdd a_43010_16058# 2.58fF
C58 CLK_IN vdd 2.08fF
C59 vbiasr vdd 33.10fF
C60 bb aa 2.62fF
C61 a_4288_11534# vdd 2.42fF
C62 a_51334_14126# a_56602_11692# 2.10fF
C63 Fvco_By4_QPH_bar vdd 2.21fF
C64 a_4226_12188# vdd 2.55fF
C65 a_50262_14152# a_51041_13108# 4.39fF
R0 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.n2 1158.04
R1 Fvco_By4_QPH_bar.t8 Fvco_By4_QPH_bar.t7 731.89
R2 Fvco_By4_QPH_bar.t3 Fvco_By4_QPH_bar.t12 719.978
R3 Fvco_By4_QPH_bar.t6 Fvco_By4_QPH_bar.t16 710.965
R4 Fvco_By4_QPH_bar.t5 Fvco_By4_QPH_bar.t17 710.965
R5 Fvco_By4_QPH_bar.t4 Fvco_By4_QPH_bar.t11 710.965
R6 Fvco_By4_QPH_bar.t16 Fvco_By4_QPH_bar.t15 579.889
R7 Fvco_By4_QPH_bar.t17 Fvco_By4_QPH_bar.t13 579.889
R8 Fvco_By4_QPH_bar.t11 Fvco_By4_QPH_bar.t10 579.889
R9 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.t5 570.03
R10 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.t4 563.963
R11 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t6 557.83
R12 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n0 458.189
R13 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.n5 435.858
R14 Fvco_By4_QPH_bar.n1 Fvco_By4_QPH_bar.t14 417.917
R15 Fvco_By4_QPH_bar.n3 Fvco_By4_QPH_bar.t9 414.213
R16 Fvco_By4_QPH_bar.n2 Fvco_By4_QPH_bar.t2 414.167
R17 Fvco_By4_QPH_bar.n6 Fvco_By4_QPH_bar.t3 245.573
R18 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.t8 244.389
R19 Fvco_By4_QPH_bar Fvco_By4_QPH_bar.n7 188.615
R20 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n4 149.023
R21 Fvco_By4_QPH_bar.n7 Fvco_By4_QPH_bar.n6 130.017
R22 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t0 69.215
R23 Fvco_By4_QPH_bar.n5 Fvco_By4_QPH_bar.n1 50.411
R24 Fvco_By4_QPH_bar.n0 Fvco_By4_QPH_bar.t1 39.949
R25 Fvco_By4_QPH_bar.n4 Fvco_By4_QPH_bar.n3 1.452
R26 a_26368_16652.t24 a_26368_16652.t50 1273.78
R27 a_26368_16652.n3 a_26368_16652.t52 182.777
R28 a_26368_16652.n3 a_26368_16652.t0 127.728
R29 a_26368_16652.t52 a_26368_16652.t21 113.753
R30 a_26368_16652.t52 a_26368_16652.t27 113.753
R31 a_26368_16652.t52 a_26368_16652.t43 113.753
R32 a_26368_16652.t52 a_26368_16652.t59 113.753
R33 a_26368_16652.t52 a_26368_16652.t53 113.753
R34 a_26368_16652.t52 a_26368_16652.t3 113.753
R35 a_26368_16652.t52 a_26368_16652.t16 113.753
R36 a_26368_16652.t52 a_26368_16652.t32 113.753
R37 a_26368_16652.t39 a_26368_16652.t28 113.753
R38 a_26368_16652.t39 a_26368_16652.t42 113.753
R39 a_26368_16652.t39 a_26368_16652.t58 113.753
R40 a_26368_16652.t39 a_26368_16652.t12 113.753
R41 a_26368_16652.n0 a_26368_16652.t35 113.753
R42 a_26368_16652.n0 a_26368_16652.t48 113.753
R43 a_26368_16652.t39 a_26368_16652.t6 113.753
R44 a_26368_16652.t39 a_26368_16652.t61 113.753
R45 a_26368_16652.t39 a_26368_16652.t13 113.753
R46 a_26368_16652.t39 a_26368_16652.t29 113.753
R47 a_26368_16652.t39 a_26368_16652.t44 113.753
R48 a_26368_16652.n0 a_26368_16652.t22 113.753
R49 a_26368_16652.n0 a_26368_16652.t54 113.753
R50 a_26368_16652.n0 a_26368_16652.t8 113.753
R51 a_26368_16652.n0 a_26368_16652.t19 113.753
R52 a_26368_16652.t39 a_26368_16652.t37 113.753
R53 a_26368_16652.t39 a_26368_16652.t33 113.753
R54 a_26368_16652.t39 a_26368_16652.t46 113.753
R55 a_26368_16652.t39 a_26368_16652.t4 113.753
R56 a_26368_16652.t39 a_26368_16652.t17 113.753
R57 a_26368_16652.n0 a_26368_16652.t36 113.753
R58 a_26368_16652.n1 a_26368_16652.t49 113.753
R59 a_26368_16652.n1 a_26368_16652.t7 113.753
R60 a_26368_16652.t39 a_26368_16652.t2 113.753
R61 a_26368_16652.t39 a_26368_16652.t14 113.753
R62 a_26368_16652.t39 a_26368_16652.t30 113.753
R63 a_26368_16652.t39 a_26368_16652.t45 113.753
R64 a_26368_16652.n0 a_26368_16652.t23 113.753
R65 a_26368_16652.n0 a_26368_16652.t55 113.753
R66 a_26368_16652.n0 a_26368_16652.t9 113.753
R67 a_26368_16652.n2 a_26368_16652.t20 113.753
R68 a_26368_16652.n2 a_26368_16652.t38 113.753
R69 a_26368_16652.n2 a_26368_16652.t34 113.753
R70 a_26368_16652.n2 a_26368_16652.t47 113.753
R71 a_26368_16652.n2 a_26368_16652.t5 113.753
R72 a_26368_16652.n2 a_26368_16652.t18 113.753
R73 a_26368_16652.t52 a_26368_16652.t51 113.753
R74 a_26368_16652.t52 a_26368_16652.t60 113.753
R75 a_26368_16652.t52 a_26368_16652.t15 113.753
R76 a_26368_16652.t52 a_26368_16652.t31 113.753
R77 a_26368_16652.t39 a_26368_16652.t26 113.753
R78 a_26368_16652.t39 a_26368_16652.t41 113.753
R79 a_26368_16652.t39 a_26368_16652.t57 113.753
R80 a_26368_16652.t39 a_26368_16652.t11 113.753
R81 a_26368_16652.t52 a_26368_16652.t56 113.753
R82 a_26368_16652.t52 a_26368_16652.t10 113.753
R83 a_26368_16652.t52 a_26368_16652.t25 113.753
R84 a_26368_16652.t52 a_26368_16652.t40 113.753
R85 a_26368_16652.t1 a_26368_16652.n3 57.482
R86 a_26368_16652.t52 a_26368_16652.n0 5.834
R87 a_26368_16652.t39 a_26368_16652.n1 3.384
R88 a_26368_16652.t52 a_26368_16652.t24 3.018
R89 a_26368_16652.t39 a_26368_16652.n2 2.785
R90 a_26368_16652.t52 a_26368_16652.t39 2.574
R91 a_23414_5032.t2 a_23414_5032.t41 1273.78
R92 a_23414_5032.n4 a_23414_5032.t14 345.988
R93 a_23414_5032.n3 a_23414_5032.t5 113.753
R94 a_23414_5032.n3 a_23414_5032.t3 113.753
R95 a_23414_5032.n3 a_23414_5032.t15 113.753
R96 a_23414_5032.n2 a_23414_5032.t36 113.753
R97 a_23414_5032.n2 a_23414_5032.t33 113.753
R98 a_23414_5032.n2 a_23414_5032.t31 113.753
R99 a_23414_5032.n2 a_23414_5032.t30 113.753
R100 a_23414_5032.n0 a_23414_5032.t7 113.753
R101 a_23414_5032.n0 a_23414_5032.t39 113.753
R102 a_23414_5032.n0 a_23414_5032.t37 113.753
R103 a_23414_5032.n0 a_23414_5032.t34 113.753
R104 a_23414_5032.n0 a_23414_5032.t45 113.753
R105 a_23414_5032.t14 a_23414_5032.t11 113.753
R106 a_23414_5032.t14 a_23414_5032.t8 113.753
R107 a_23414_5032.t14 a_23414_5032.t6 113.753
R108 a_23414_5032.t14 a_23414_5032.t4 113.753
R109 a_23414_5032.n0 a_23414_5032.t21 113.753
R110 a_23414_5032.n0 a_23414_5032.t17 113.753
R111 a_23414_5032.n1 a_23414_5032.t35 113.753
R112 a_23414_5032.n1 a_23414_5032.t56 113.753
R113 a_23414_5032.n1 a_23414_5032.t51 113.753
R114 a_23414_5032.n1 a_23414_5032.t49 113.753
R115 a_23414_5032.n1 a_23414_5032.t47 113.753
R116 a_23414_5032.n0 a_23414_5032.t24 113.753
R117 a_23414_5032.n0 a_23414_5032.t58 113.753
R118 a_23414_5032.n0 a_23414_5032.t55 113.753
R119 a_23414_5032.n0 a_23414_5032.t52 113.753
R120 a_23414_5032.t14 a_23414_5032.t9 113.753
R121 a_23414_5032.t14 a_23414_5032.t28 113.753
R122 a_23414_5032.t14 a_23414_5032.t25 113.753
R123 a_23414_5032.t14 a_23414_5032.t23 113.753
R124 a_23414_5032.t14 a_23414_5032.t20 113.753
R125 a_23414_5032.n0 a_23414_5032.t27 113.753
R126 a_23414_5032.t14 a_23414_5032.t26 113.753
R127 a_23414_5032.t14 a_23414_5032.t42 113.753
R128 a_23414_5032.t14 a_23414_5032.t60 113.753
R129 a_23414_5032.t14 a_23414_5032.t59 113.753
R130 a_23414_5032.t14 a_23414_5032.t57 113.753
R131 a_23414_5032.t14 a_23414_5032.t54 113.753
R132 a_23414_5032.n0 a_23414_5032.t29 113.753
R133 a_23414_5032.n0 a_23414_5032.t13 113.753
R134 a_23414_5032.n0 a_23414_5032.t12 113.753
R135 a_23414_5032.t14 a_23414_5032.t10 113.753
R136 a_23414_5032.t14 a_23414_5032.t19 113.753
R137 a_23414_5032.t14 a_23414_5032.t44 113.753
R138 a_23414_5032.t14 a_23414_5032.t43 113.753
R139 a_23414_5032.t14 a_23414_5032.t40 113.753
R140 a_23414_5032.t14 a_23414_5032.t38 113.753
R141 a_23414_5032.n0 a_23414_5032.t22 113.753
R142 a_23414_5032.n0 a_23414_5032.t18 113.753
R143 a_23414_5032.n0 a_23414_5032.t16 113.753
R144 a_23414_5032.t14 a_23414_5032.t32 113.753
R145 a_23414_5032.t14 a_23414_5032.t53 113.753
R146 a_23414_5032.t14 a_23414_5032.t50 113.753
R147 a_23414_5032.t14 a_23414_5032.t48 113.753
R148 a_23414_5032.t14 a_23414_5032.t46 113.753
R149 a_23414_5032.t0 a_23414_5032.n5 82.513
R150 a_23414_5032.n4 a_23414_5032.t1 28.697
R151 a_23414_5032.t14 a_23414_5032.n0 4.31
R152 a_23414_5032.n5 a_23414_5032.n4 3.507
R153 a_23414_5032.n0 a_23414_5032.n3 3.224
R154 a_23414_5032.t14 a_23414_5032.n1 2.869
R155 a_23414_5032.t14 a_23414_5032.n2 2.708
R156 a_23414_5032.n5 a_23414_5032.t2 2.634
R157 a_26690_784.n1 a_26690_784.t2 434.481
R158 a_26690_784.n0 a_26690_784.t3 217.163
R159 a_26690_784.t1 a_26690_784.n1 52.152
R160 a_26690_784.n0 a_26690_784.t0 3.106
R161 a_26690_784.n1 a_26690_784.n0 0.879
R162 vinit.n15 vinit.n14 70.035
R163 vinit.n9 vinit.t44 56.95
R164 vinit.n11 vinit.t42 56.876
R165 vinit.n12 vinit.t43 56.876
R166 vinit.n10 vinit.t40 56.876
R167 vinit.n9 vinit.t41 56.876
R168 vinit.n15 vinit.t30 7.425
R169 vinit.n34 vinit.t21 7.425
R170 vinit.n32 vinit.t25 5.713
R171 vinit.n32 vinit.t31 5.713
R172 vinit.n30 vinit.t29 5.713
R173 vinit.n30 vinit.t34 5.713
R174 vinit.n28 vinit.t37 5.713
R175 vinit.n28 vinit.t23 5.713
R176 vinit.n26 vinit.t28 5.713
R177 vinit.n26 vinit.t27 5.713
R178 vinit.n24 vinit.t33 5.713
R179 vinit.n24 vinit.t36 5.713
R180 vinit.n22 vinit.t22 5.713
R181 vinit.n22 vinit.t20 5.713
R182 vinit.n20 vinit.t26 5.713
R183 vinit.n20 vinit.t32 5.713
R184 vinit.n16 vinit.t38 5.713
R185 vinit.n16 vinit.t24 5.713
R186 vinit.n18 vinit.t35 5.713
R187 vinit.n18 vinit.t39 5.713
R188 vinit.n45 vinit.t17 5.244
R189 vinit.n35 vinit.t0 5.244
R190 vinit.n0 vinit.t14 3.48
R191 vinit.n0 vinit.t1 3.48
R192 vinit.n1 vinit.t6 3.48
R193 vinit.n1 vinit.t5 3.48
R194 vinit.n2 vinit.t13 3.48
R195 vinit.n2 vinit.t11 3.48
R196 vinit.n3 vinit.t19 3.48
R197 vinit.n3 vinit.t4 3.48
R198 vinit.n4 vinit.t3 3.48
R199 vinit.n4 vinit.t10 3.48
R200 vinit.n5 vinit.t9 3.48
R201 vinit.n5 vinit.t18 3.48
R202 vinit.n6 vinit.t16 3.48
R203 vinit.n6 vinit.t2 3.48
R204 vinit.n7 vinit.t8 3.48
R205 vinit.n7 vinit.t7 3.48
R206 vinit.n8 vinit.t15 3.48
R207 vinit.n8 vinit.t12 3.48
R208 vinit.n41 vinit.n3 1.766
R209 vinit.n44 vinit.n0 1.766
R210 vinit.n38 vinit.n6 1.766
R211 vinit.n37 vinit.n7 1.764
R212 vinit.n40 vinit.n4 1.762
R213 vinit.n42 vinit.n2 1.761
R214 vinit.n39 vinit.n5 1.758
R215 vinit.n43 vinit.n1 1.758
R216 vinit.n36 vinit.n8 1.754
R217 vinit.n23 vinit.n22 1.714
R218 vinit.n17 vinit.n16 1.714
R219 vinit.n29 vinit.n28 1.714
R220 vinit.n31 vinit.n30 1.712
R221 vinit.n25 vinit.n24 1.71
R222 vinit.n21 vinit.n20 1.709
R223 vinit.n27 vinit.n26 1.706
R224 vinit.n19 vinit.n18 1.706
R225 vinit.n33 vinit.n32 1.702
R226 vinit vinit.n45 0.543
R227 vinit.n14 vinit.n13 0.322
R228 vinit.n35 vinit.n34 0.295
R229 vinit.n12 vinit.n11 0.073
R230 vinit.n10 vinit.n9 0.073
R231 vinit.n13 vinit.n12 0.051
R232 vinit.n34 vinit.n33 0.032
R233 vinit.n40 vinit.n39 0.031
R234 vinit.n27 vinit.n25 0.031
R235 vinit.n43 vinit.n42 0.031
R236 vinit.n21 vinit.n19 0.031
R237 vinit.n37 vinit.n36 0.031
R238 vinit.n33 vinit.n31 0.031
R239 vinit.n36 vinit.n35 0.031
R240 vinit.n44 vinit.n43 0.03
R241 vinit.n19 vinit.n17 0.03
R242 vinit.n45 vinit.n44 0.03
R243 vinit.n17 vinit.n15 0.03
R244 vinit.n38 vinit.n37 0.03
R245 vinit.n31 vinit.n29 0.03
R246 vinit.n41 vinit.n40 0.03
R247 vinit.n25 vinit.n23 0.03
R248 vinit.n42 vinit.n41 0.03
R249 vinit.n23 vinit.n21 0.03
R250 vinit.n39 vinit.n38 0.03
R251 vinit.n29 vinit.n27 0.03
R252 vinit.n13 vinit.n10 0.022
R253 a_14188_14050.t12 a_14188_14050.t53 1273.78
R254 a_14188_14050.n3 a_14188_14050.t31 161.992
R255 a_14188_14050.t39 a_14188_14050.t40 113.753
R256 a_14188_14050.t39 a_14188_14050.t50 113.753
R257 a_14188_14050.t39 a_14188_14050.t47 113.753
R258 a_14188_14050.t39 a_14188_14050.t11 113.753
R259 a_14188_14050.n0 a_14188_14050.t23 113.753
R260 a_14188_14050.n0 a_14188_14050.t6 113.753
R261 a_14188_14050.n0 a_14188_14050.t19 113.753
R262 a_14188_14050.n0 a_14188_14050.t41 113.753
R263 a_14188_14050.t39 a_14188_14050.t55 113.753
R264 a_14188_14050.t39 a_14188_14050.t9 113.753
R265 a_14188_14050.t39 a_14188_14050.t8 113.753
R266 a_14188_14050.t39 a_14188_14050.t26 113.753
R267 a_14188_14050.n0 a_14188_14050.t42 113.753
R268 a_14188_14050.n0 a_14188_14050.t24 113.753
R269 a_14188_14050.n0 a_14188_14050.t38 113.753
R270 a_14188_14050.n0 a_14188_14050.t57 113.753
R271 a_14188_14050.t31 a_14188_14050.t21 113.753
R272 a_14188_14050.t31 a_14188_14050.t36 113.753
R273 a_14188_14050.t31 a_14188_14050.t33 113.753
R274 a_14188_14050.t31 a_14188_14050.t56 113.753
R275 a_14188_14050.n0 a_14188_14050.t10 113.753
R276 a_14188_14050.n0 a_14188_14050.t51 113.753
R277 a_14188_14050.n0 a_14188_14050.t5 113.753
R278 a_14188_14050.n0 a_14188_14050.t25 113.753
R279 a_14188_14050.t31 a_14188_14050.t49 113.753
R280 a_14188_14050.t31 a_14188_14050.t4 113.753
R281 a_14188_14050.t31 a_14188_14050.t60 113.753
R282 a_14188_14050.t31 a_14188_14050.t22 113.753
R283 a_14188_14050.n1 a_14188_14050.t37 113.753
R284 a_14188_14050.n1 a_14188_14050.t18 113.753
R285 a_14188_14050.n1 a_14188_14050.t30 113.753
R286 a_14188_14050.n1 a_14188_14050.t54 113.753
R287 a_14188_14050.n2 a_14188_14050.t3 113.753
R288 a_14188_14050.n2 a_14188_14050.t16 113.753
R289 a_14188_14050.n2 a_14188_14050.t14 113.753
R290 a_14188_14050.n2 a_14188_14050.t35 113.753
R291 a_14188_14050.n0 a_14188_14050.t48 113.753
R292 a_14188_14050.n0 a_14188_14050.t29 113.753
R293 a_14188_14050.n0 a_14188_14050.t45 113.753
R294 a_14188_14050.n0 a_14188_14050.t7 113.753
R295 a_14188_14050.t31 a_14188_14050.t46 113.753
R296 a_14188_14050.t31 a_14188_14050.t61 113.753
R297 a_14188_14050.t31 a_14188_14050.t59 113.753
R298 a_14188_14050.t31 a_14188_14050.t20 113.753
R299 a_14188_14050.t31 a_14188_14050.t28 113.753
R300 a_14188_14050.t31 a_14188_14050.t44 113.753
R301 a_14188_14050.t31 a_14188_14050.t43 113.753
R302 a_14188_14050.t31 a_14188_14050.t2 113.753
R303 a_14188_14050.n0 a_14188_14050.t15 113.753
R304 a_14188_14050.n0 a_14188_14050.t58 113.753
R305 a_14188_14050.n0 a_14188_14050.t13 113.753
R306 a_14188_14050.n0 a_14188_14050.t32 113.753
R307 a_14188_14050.t31 a_14188_14050.t34 113.753
R308 a_14188_14050.t31 a_14188_14050.t17 113.753
R309 a_14188_14050.t31 a_14188_14050.t27 113.753
R310 a_14188_14050.n0 a_14188_14050.t52 113.753
R311 a_14188_14050.t1 a_14188_14050.n4 57.821
R312 a_14188_14050.n3 a_14188_14050.t0 47.07
R313 a_14188_14050.n4 a_14188_14050.t12 6.878
R314 a_14188_14050.n4 a_14188_14050.n3 3.96
R315 a_14188_14050.t31 a_14188_14050.t39 3.88
R316 a_14188_14050.t31 a_14188_14050.n0 3.25
R317 a_14188_14050.n0 a_14188_14050.n1 2.856
R318 a_14188_14050.t31 a_14188_14050.n2 2.454
R319 a_49874_4150.n0 a_49874_4150.t12 19.742
R320 a_49874_4150.n0 a_49874_4150.t6 18.733
R321 a_49874_4150.t3 a_49874_4150.n1 18.498
R322 a_49874_4150.n3 a_49874_4150.t2 17.928
R323 a_49874_4150.n0 a_49874_4150.t9 16.208
R324 a_49874_4150.n1 a_49874_4150.t1 15.946
R325 a_49874_4150.n2 a_49874_4150.t5 9.424
R326 a_49874_4150.n2 a_49874_4150.t8 8.34
R327 a_49874_4150.n2 a_49874_4150.t11 5.724
R328 a_49874_4150.n1 a_49874_4150.t0 5.514
R329 a_49874_4150.n0 a_49874_4150.t4 5.514
R330 a_49874_4150.n3 a_49874_4150.t7 5.512
R331 a_49874_4150.n1 a_49874_4150.n0 4.479
R332 a_49874_4150.n4 a_49874_4150.n3 4.094
R333 a_49874_4150.n4 a_49874_4150.t10 3.856
R334 a_49874_4150.n0 a_49874_4150.n4 3.301
R335 a_49874_4150.n0 a_49874_4150.n2 2.294
R336 Fvco_By4_QPH.t10 Fvco_By4_QPH.t19 731.89
R337 Fvco_By4_QPH.t14 Fvco_By4_QPH.t6 731.89
R338 Fvco_By4_QPH.t3 Fvco_By4_QPH.t13 731.89
R339 Fvco_By4_QPH.t5 Fvco_By4_QPH.t16 718.506
R340 Fvco_By4_QPH.t11 Fvco_By4_QPH.t15 710.965
R341 Fvco_By4_QPH.t7 Fvco_By4_QPH.t14 622.637
R342 Fvco_By4_QPH.n8 Fvco_By4_QPH.n7 617.524
R343 Fvco_By4_QPH.n4 Fvco_By4_QPH.n3 580.872
R344 Fvco_By4_QPH.t15 Fvco_By4_QPH.t2 579.889
R345 Fvco_By4_QPH.n3 Fvco_By4_QPH.t12 491.229
R346 Fvco_By4_QPH.n4 Fvco_By4_QPH.t4 489.182
R347 Fvco_By4_QPH.n9 Fvco_By4_QPH.t11 418.965
R348 Fvco_By4_QPH.n8 Fvco_By4_QPH.t18 414.13
R349 Fvco_By4_QPH.n5 Fvco_By4_QPH.t9 349.273
R350 Fvco_By4_QPH.n2 Fvco_By4_QPH.t8 333.651
R351 Fvco_By4_QPH.n6 Fvco_By4_QPH.t3 317.894
R352 Fvco_By4_QPH.n2 Fvco_By4_QPH.t17 297.233
R353 Fvco_By4_QPH.n6 Fvco_By4_QPH.t5 291.323
R354 Fvco_By4_QPH.n5 Fvco_By4_QPH.t10 252.624
R355 Fvco_By4_QPH.n3 Fvco_By4_QPH.t7 227.612
R356 Fvco_By4_QPH.t9 Fvco_By4_QPH.n4 227.612
R357 Fvco_By4_QPH.n7 Fvco_By4_QPH.n5 198.896
R358 Fvco_By4_QPH.n9 Fvco_By4_QPH.n8 152.778
R359 Fvco_By4_QPH.n0 Fvco_By4_QPH.t1 92.046
R360 Fvco_By4_QPH.n1 Fvco_By4_QPH.n2 70.221
R361 Fvco_By4_QPH.n0 Fvco_By4_QPH.t0 61.427
R362 Fvco_By4_QPH Fvco_By4_QPH.n9 38.508
R363 Fvco_By4_QPH.n7 Fvco_By4_QPH.n6 31.687
R364 Fvco_By4_QPH Fvco_By4_QPH.n1 10.972
R365 Fvco_By4_QPH.n1 Fvco_By4_QPH.n0 0.154
R366 a_26036_4988.t16 a_26036_4988.t22 1273.78
R367 a_26036_4988.n0 a_26036_4988.t44 415.476
R368 a_26036_4988.t44 a_26036_4988.t37 113.753
R369 a_26036_4988.t44 a_26036_4988.t34 113.753
R370 a_26036_4988.t44 a_26036_4988.t32 113.753
R371 a_26036_4988.t20 a_26036_4988.t46 113.753
R372 a_26036_4988.t20 a_26036_4988.t7 113.753
R373 a_26036_4988.t20 a_26036_4988.t4 113.753
R374 a_26036_4988.t20 a_26036_4988.t61 113.753
R375 a_26036_4988.t44 a_26036_4988.t14 113.753
R376 a_26036_4988.t44 a_26036_4988.t47 113.753
R377 a_26036_4988.t44 a_26036_4988.t10 113.753
R378 a_26036_4988.t44 a_26036_4988.t6 113.753
R379 a_26036_4988.t44 a_26036_4988.t3 113.753
R380 a_26036_4988.t20 a_26036_4988.t15 113.753
R381 a_26036_4988.t20 a_26036_4988.t41 113.753
R382 a_26036_4988.t20 a_26036_4988.t38 113.753
R383 a_26036_4988.t20 a_26036_4988.t35 113.753
R384 a_26036_4988.n1 a_26036_4988.t55 113.753
R385 a_26036_4988.n1 a_26036_4988.t52 113.753
R386 a_26036_4988.t20 a_26036_4988.t49 113.753
R387 a_26036_4988.t20 a_26036_4988.t5 113.753
R388 a_26036_4988.t20 a_26036_4988.t27 113.753
R389 a_26036_4988.t20 a_26036_4988.t25 113.753
R390 a_26036_4988.t20 a_26036_4988.t18 113.753
R391 a_26036_4988.n1 a_26036_4988.t36 113.753
R392 a_26036_4988.n1 a_26036_4988.t8 113.753
R393 a_26036_4988.n1 a_26036_4988.t29 113.753
R394 a_26036_4988.n1 a_26036_4988.t26 113.753
R395 a_26036_4988.t20 a_26036_4988.t23 113.753
R396 a_26036_4988.t20 a_26036_4988.t39 113.753
R397 a_26036_4988.t20 a_26036_4988.t59 113.753
R398 a_26036_4988.t20 a_26036_4988.t57 113.753
R399 a_26036_4988.t20 a_26036_4988.t53 113.753
R400 a_26036_4988.n1 a_26036_4988.t60 113.753
R401 a_26036_4988.t20 a_26036_4988.t58 113.753
R402 a_26036_4988.t20 a_26036_4988.t56 113.753
R403 a_26036_4988.t20 a_26036_4988.t11 113.753
R404 a_26036_4988.t20 a_26036_4988.t31 113.753
R405 a_26036_4988.t20 a_26036_4988.t30 113.753
R406 a_26036_4988.t20 a_26036_4988.t28 113.753
R407 a_26036_4988.n1 a_26036_4988.t42 113.753
R408 a_26036_4988.n1 a_26036_4988.t19 113.753
R409 a_26036_4988.n1 a_26036_4988.t45 113.753
R410 a_26036_4988.n2 a_26036_4988.t43 113.753
R411 a_26036_4988.n2 a_26036_4988.t40 113.753
R412 a_26036_4988.n2 a_26036_4988.t51 113.753
R413 a_26036_4988.n2 a_26036_4988.t13 113.753
R414 a_26036_4988.n2 a_26036_4988.t12 113.753
R415 a_26036_4988.n2 a_26036_4988.t9 113.753
R416 a_26036_4988.t44 a_26036_4988.t33 113.753
R417 a_26036_4988.t44 a_26036_4988.t54 113.753
R418 a_26036_4988.t44 a_26036_4988.t50 113.753
R419 a_26036_4988.t44 a_26036_4988.t48 113.753
R420 a_26036_4988.t44 a_26036_4988.t2 113.753
R421 a_26036_4988.t44 a_26036_4988.t24 113.753
R422 a_26036_4988.t44 a_26036_4988.t21 113.753
R423 a_26036_4988.t44 a_26036_4988.t17 113.753
R424 a_26036_4988.t1 a_26036_4988.n0 81.094
R425 a_26036_4988.n0 a_26036_4988.t0 28.577
R426 a_26036_4988.t44 a_26036_4988.n1 6.49
R427 a_26036_4988.n0 a_26036_4988.t16 5.37
R428 a_26036_4988.t20 a_26036_4988.n2 4.699
R429 a_26036_4988.t44 a_26036_4988.t20 2.967
R430 a_25099_11445.t53 a_25099_11445.t41 1273.78
R431 a_25099_11445.n3 a_25099_11445.t40 218.051
R432 a_25099_11445.t40 a_25099_11445.t49 113.753
R433 a_25099_11445.t40 a_25099_11445.t8 113.753
R434 a_25099_11445.t40 a_25099_11445.t29 113.753
R435 a_25099_11445.t40 a_25099_11445.t21 113.753
R436 a_25099_11445.t40 a_25099_11445.t42 113.753
R437 a_25099_11445.t40 a_25099_11445.t59 113.753
R438 a_25099_11445.t40 a_25099_11445.t57 113.753
R439 a_25099_11445.n2 a_25099_11445.t6 113.753
R440 a_25099_11445.n2 a_25099_11445.t16 113.753
R441 a_25099_11445.n2 a_25099_11445.t37 113.753
R442 a_25099_11445.n2 a_25099_11445.t54 113.753
R443 a_25099_11445.t40 a_25099_11445.t19 113.753
R444 a_25099_11445.n0 a_25099_11445.t51 113.753
R445 a_25099_11445.n0 a_25099_11445.t10 113.753
R446 a_25099_11445.n0 a_25099_11445.t31 113.753
R447 a_25099_11445.n1 a_25099_11445.t26 113.753
R448 a_25099_11445.n1 a_25099_11445.t35 113.753
R449 a_25099_11445.n1 a_25099_11445.t47 113.753
R450 a_25099_11445.n1 a_25099_11445.t4 113.753
R451 a_25099_11445.n1 a_25099_11445.t23 113.753
R452 a_25099_11445.n0 a_25099_11445.t43 113.753
R453 a_25099_11445.n0 a_25099_11445.t60 113.753
R454 a_25099_11445.t15 a_25099_11445.t58 113.753
R455 a_25099_11445.t15 a_25099_11445.t7 113.753
R456 a_25099_11445.t15 a_25099_11445.t17 113.753
R457 a_25099_11445.t15 a_25099_11445.t38 113.753
R458 a_25099_11445.t15 a_25099_11445.t55 113.753
R459 a_25099_11445.n0 a_25099_11445.t20 113.753
R460 a_25099_11445.n0 a_25099_11445.t52 113.753
R461 a_25099_11445.n0 a_25099_11445.t11 113.753
R462 a_25099_11445.t15 a_25099_11445.t32 113.753
R463 a_25099_11445.t15 a_25099_11445.t27 113.753
R464 a_25099_11445.t15 a_25099_11445.t36 113.753
R465 a_25099_11445.t15 a_25099_11445.t48 113.753
R466 a_25099_11445.t15 a_25099_11445.t5 113.753
R467 a_25099_11445.t15 a_25099_11445.t24 113.753
R468 a_25099_11445.t15 a_25099_11445.t39 113.753
R469 a_25099_11445.t15 a_25099_11445.t56 113.753
R470 a_25099_11445.t15 a_25099_11445.t12 113.753
R471 a_25099_11445.n0 a_25099_11445.t44 113.753
R472 a_25099_11445.n0 a_25099_11445.t61 113.753
R473 a_25099_11445.t15 a_25099_11445.t14 113.753
R474 a_25099_11445.t15 a_25099_11445.t13 113.753
R475 a_25099_11445.t15 a_25099_11445.t28 113.753
R476 a_25099_11445.t40 a_25099_11445.t50 113.753
R477 a_25099_11445.t40 a_25099_11445.t9 113.753
R478 a_25099_11445.t40 a_25099_11445.t30 113.753
R479 a_25099_11445.t40 a_25099_11445.t25 113.753
R480 a_25099_11445.t15 a_25099_11445.t34 113.753
R481 a_25099_11445.t15 a_25099_11445.t46 113.753
R482 a_25099_11445.t15 a_25099_11445.t3 113.753
R483 a_25099_11445.t15 a_25099_11445.t22 113.753
R484 a_25099_11445.t40 a_25099_11445.t33 113.753
R485 a_25099_11445.t40 a_25099_11445.t45 113.753
R486 a_25099_11445.t40 a_25099_11445.t2 113.753
R487 a_25099_11445.t40 a_25099_11445.t18 113.753
R488 a_25099_11445.t0 a_25099_11445.n4 56.779
R489 a_25099_11445.n3 a_25099_11445.t1 28.581
R490 a_25099_11445.t40 a_25099_11445.n0 5.834
R491 a_25099_11445.n4 a_25099_11445.t53 4.799
R492 a_25099_11445.n4 a_25099_11445.n3 3.709
R493 a_25099_11445.t15 a_25099_11445.n1 2.869
R494 a_25099_11445.t40 a_25099_11445.t15 2.816
R495 a_25099_11445.t15 a_25099_11445.n2 2.586
R496 a_17685_3840.n28 a_17685_3840.n27 660.793
R497 a_17685_3840.n58 a_17685_3840.n57 649.743
R498 a_17685_3840.n61 a_17685_3840.n60 574.593
R499 a_17685_3840.n29 a_17685_3840.n28 416.406
R500 a_17685_3840.n62 a_17685_3840.n61 415.789
R501 a_17685_3840.n25 a_17685_3840.n24 270.636
R502 a_17685_3840.n27 a_17685_3840.n26 262.3
R503 a_17685_3840.n28 a_17685_3840.n25 198.935
R504 a_17685_3840.n60 a_17685_3840.t12 197.212
R505 a_17685_3840.n26 a_17685_3840.t6 185.816
R506 a_17685_3840.n27 a_17685_3840.t16 176.327
R507 a_17685_3840.n59 a_17685_3840.t11 173.989
R508 a_17685_3840.n25 a_17685_3840.t13 154.605
R509 a_17685_3840.n24 a_17685_3840.t14 151.674
R510 a_17685_3840.n63 a_17685_3840.t15 118.032
R511 a_17685_3840.n61 a_17685_3840.n59 107.97
R512 a_17685_3840.n30 a_17685_3840.n29 104.297
R513 a_17685_3840.n64 a_17685_3840.n63 103.649
R514 a_17685_3840.n68 a_17685_3840.n67 100.879
R515 a_17685_3840.n65 a_17685_3840.n64 83.404
R516 a_17685_3840.n65 a_17685_3840.t5 81.437
R517 a_17685_3840.n30 a_17685_3840.t10 69.653
R518 a_17685_3840.n31 a_17685_3840.t2 68.683
R519 a_17685_3840.n64 a_17685_3840.n34 66.545
R520 a_17685_3840.n63 a_17685_3840.n62 47.861
R521 a_17685_3840.n23 a_17685_3840.n22 45.936
R522 a_17685_3840.n31 a_17685_3840.n30 45.7
R523 a_17685_3840.n29 a_17685_3840.n23 41.108
R524 a_17685_3840.n62 a_17685_3840.n58 41.07
R525 a_17685_3840.n66 a_17685_3840.n32 40.118
R526 a_17685_3840.n34 a_17685_3840.t9 28.576
R527 a_17685_3840.n33 a_17685_3840.t7 28.565
R528 a_17685_3840.n33 a_17685_3840.t8 28.565
R529 a_17685_3840.n32 a_17685_3840.t3 28.565
R530 a_17685_3840.n32 a_17685_3840.t0 28.565
R531 a_17685_3840.n68 a_17685_3840.t1 28.565
R532 a_17685_3840.t4 a_17685_3840.n68 28.565
R533 a_17685_3840.n57 a_17685_3840.n45 24.999
R534 a_17685_3840.n66 a_17685_3840.n65 24.605
R535 a_17685_3840.n22 a_17685_3840.n10 24.399
R536 a_17685_3840.n35 a_17685_3840.t50 23.529
R537 a_17685_3840.n0 a_17685_3840.t43 23.485
R538 a_17685_3840.n11 a_17685_3840.t35 23.474
R539 a_17685_3840.n46 a_17685_3840.t59 23.456
R540 a_17685_3840.n67 a_17685_3840.n66 20.217
R541 a_17685_3840.n67 a_17685_3840.n31 19.791
R542 a_17685_3840.n45 a_17685_3840.t39 15.401
R543 a_17685_3840.n10 a_17685_3840.t54 15.374
R544 a_17685_3840.n56 a_17685_3840.t26 15.341
R545 a_17685_3840.n21 a_17685_3840.t27 15.334
R546 a_17685_3840.n22 a_17685_3840.n21 12.228
R547 a_17685_3840.n57 a_17685_3840.n56 11.433
R548 a_17685_3840.n44 a_17685_3840.n43 10.674
R549 a_17685_3840.n43 a_17685_3840.n42 10.674
R550 a_17685_3840.n42 a_17685_3840.n41 10.674
R551 a_17685_3840.n41 a_17685_3840.n40 10.674
R552 a_17685_3840.n40 a_17685_3840.n39 10.674
R553 a_17685_3840.n39 a_17685_3840.n38 10.674
R554 a_17685_3840.n38 a_17685_3840.n37 10.674
R555 a_17685_3840.n37 a_17685_3840.n36 10.674
R556 a_17685_3840.n36 a_17685_3840.n35 10.674
R557 a_17685_3840.n20 a_17685_3840.n19 10.655
R558 a_17685_3840.n19 a_17685_3840.n18 10.655
R559 a_17685_3840.n18 a_17685_3840.n17 10.655
R560 a_17685_3840.n17 a_17685_3840.n16 10.655
R561 a_17685_3840.n16 a_17685_3840.n15 10.655
R562 a_17685_3840.n15 a_17685_3840.n14 10.655
R563 a_17685_3840.n14 a_17685_3840.n13 10.655
R564 a_17685_3840.n13 a_17685_3840.n12 10.655
R565 a_17685_3840.n12 a_17685_3840.n11 10.655
R566 a_17685_3840.n9 a_17685_3840.n8 10.637
R567 a_17685_3840.n8 a_17685_3840.n7 10.637
R568 a_17685_3840.n7 a_17685_3840.n6 10.637
R569 a_17685_3840.n6 a_17685_3840.n5 10.637
R570 a_17685_3840.n5 a_17685_3840.n4 10.637
R571 a_17685_3840.n4 a_17685_3840.n3 10.637
R572 a_17685_3840.n3 a_17685_3840.n2 10.637
R573 a_17685_3840.n2 a_17685_3840.n1 10.637
R574 a_17685_3840.n1 a_17685_3840.n0 10.637
R575 a_17685_3840.n55 a_17685_3840.n54 10.625
R576 a_17685_3840.n54 a_17685_3840.n53 10.625
R577 a_17685_3840.n53 a_17685_3840.n52 10.625
R578 a_17685_3840.n52 a_17685_3840.n51 10.625
R579 a_17685_3840.n51 a_17685_3840.n50 10.625
R580 a_17685_3840.n50 a_17685_3840.n49 10.625
R581 a_17685_3840.n49 a_17685_3840.n48 10.625
R582 a_17685_3840.n48 a_17685_3840.n47 10.625
R583 a_17685_3840.n47 a_17685_3840.n46 10.625
R584 a_17685_3840.n46 a_17685_3840.t19 8.716
R585 a_17685_3840.n47 a_17685_3840.t25 8.716
R586 a_17685_3840.n48 a_17685_3840.t34 8.716
R587 a_17685_3840.n49 a_17685_3840.t40 8.716
R588 a_17685_3840.n50 a_17685_3840.t17 8.716
R589 a_17685_3840.n51 a_17685_3840.t23 8.716
R590 a_17685_3840.n52 a_17685_3840.t32 8.716
R591 a_17685_3840.n53 a_17685_3840.t30 8.716
R592 a_17685_3840.n54 a_17685_3840.t37 8.716
R593 a_17685_3840.n55 a_17685_3840.t45 8.716
R594 a_17685_3840.n0 a_17685_3840.t51 8.713
R595 a_17685_3840.n1 a_17685_3840.t56 8.713
R596 a_17685_3840.n2 a_17685_3840.t64 8.713
R597 a_17685_3840.n3 a_17685_3840.t20 8.713
R598 a_17685_3840.n4 a_17685_3840.t48 8.713
R599 a_17685_3840.n5 a_17685_3840.t53 8.713
R600 a_17685_3840.n6 a_17685_3840.t60 8.713
R601 a_17685_3840.n7 a_17685_3840.t58 8.713
R602 a_17685_3840.n8 a_17685_3840.t63 8.713
R603 a_17685_3840.n9 a_17685_3840.t22 8.713
R604 a_17685_3840.n11 a_17685_3840.t42 8.708
R605 a_17685_3840.n12 a_17685_3840.t49 8.708
R606 a_17685_3840.n13 a_17685_3840.t55 8.708
R607 a_17685_3840.n14 a_17685_3840.t61 8.708
R608 a_17685_3840.n15 a_17685_3840.t18 8.708
R609 a_17685_3840.n16 a_17685_3840.t24 8.708
R610 a_17685_3840.n17 a_17685_3840.t33 8.708
R611 a_17685_3840.n18 a_17685_3840.t31 8.708
R612 a_17685_3840.n19 a_17685_3840.t38 8.708
R613 a_17685_3840.n20 a_17685_3840.t46 8.708
R614 a_17685_3840.n44 a_17685_3840.t52 8.704
R615 a_17685_3840.n35 a_17685_3840.t57 8.704
R616 a_17685_3840.n36 a_17685_3840.t62 8.704
R617 a_17685_3840.n37 a_17685_3840.t21 8.704
R618 a_17685_3840.n38 a_17685_3840.t28 8.704
R619 a_17685_3840.n39 a_17685_3840.t29 8.704
R620 a_17685_3840.n40 a_17685_3840.t36 8.704
R621 a_17685_3840.n41 a_17685_3840.t44 8.704
R622 a_17685_3840.n42 a_17685_3840.t41 8.704
R623 a_17685_3840.n43 a_17685_3840.t47 8.704
R624 a_17685_3840.n21 a_17685_3840.n20 8.14
R625 a_17685_3840.n45 a_17685_3840.n44 8.128
R626 a_17685_3840.n56 a_17685_3840.n55 8.116
R627 a_17685_3840.n10 a_17685_3840.n9 8.112
R628 a_17685_3840.n34 a_17685_3840.n33 0.712
R629 a_14266_8900.t16 a_14266_8900.t25 1273.78
R630 a_14266_8900.n3 a_14266_8900.t54 193.916
R631 a_14266_8900.t54 a_14266_8900.t21 113.753
R632 a_14266_8900.t54 a_14266_8900.t11 113.753
R633 a_14266_8900.t54 a_14266_8900.t32 113.753
R634 a_14266_8900.t54 a_14266_8900.t41 113.753
R635 a_14266_8900.t54 a_14266_8900.t52 113.753
R636 a_14266_8900.t54 a_14266_8900.t50 113.753
R637 a_14266_8900.t54 a_14266_8900.t59 113.753
R638 a_14266_8900.t54 a_14266_8900.t18 113.753
R639 a_14266_8900.n2 a_14266_8900.t8 113.753
R640 a_14266_8900.n2 a_14266_8900.t48 113.753
R641 a_14266_8900.n2 a_14266_8900.t42 113.753
R642 a_14266_8900.n2 a_14266_8900.t55 113.753
R643 a_14266_8900.n0 a_14266_8900.t17 113.753
R644 a_14266_8900.n0 a_14266_8900.t34 113.753
R645 a_14266_8900.n1 a_14266_8900.t45 113.753
R646 a_14266_8900.n1 a_14266_8900.t39 113.753
R647 a_14266_8900.n1 a_14266_8900.t13 113.753
R648 a_14266_8900.n1 a_14266_8900.t5 113.753
R649 a_14266_8900.n1 a_14266_8900.t29 113.753
R650 a_14266_8900.n0 a_14266_8900.t23 113.753
R651 a_14266_8900.n0 a_14266_8900.t53 113.753
R652 a_14266_8900.n0 a_14266_8900.t51 113.753
R653 a_14266_8900.n0 a_14266_8900.t60 113.753
R654 a_14266_8900.t47 a_14266_8900.t20 113.753
R655 a_14266_8900.t47 a_14266_8900.t9 113.753
R656 a_14266_8900.t47 a_14266_8900.t49 113.753
R657 a_14266_8900.t47 a_14266_8900.t43 113.753
R658 a_14266_8900.t47 a_14266_8900.t56 113.753
R659 a_14266_8900.n0 a_14266_8900.t19 113.753
R660 a_14266_8900.t47 a_14266_8900.t35 113.753
R661 a_14266_8900.t47 a_14266_8900.t46 113.753
R662 a_14266_8900.t47 a_14266_8900.t40 113.753
R663 a_14266_8900.t47 a_14266_8900.t14 113.753
R664 a_14266_8900.t47 a_14266_8900.t6 113.753
R665 a_14266_8900.t47 a_14266_8900.t30 113.753
R666 a_14266_8900.n0 a_14266_8900.t24 113.753
R667 a_14266_8900.n0 a_14266_8900.t2 113.753
R668 a_14266_8900.n0 a_14266_8900.t61 113.753
R669 a_14266_8900.t47 a_14266_8900.t27 113.753
R670 a_14266_8900.t47 a_14266_8900.t36 113.753
R671 a_14266_8900.t47 a_14266_8900.t31 113.753
R672 a_14266_8900.t47 a_14266_8900.t58 113.753
R673 a_14266_8900.t47 a_14266_8900.t57 113.753
R674 a_14266_8900.t47 a_14266_8900.t7 113.753
R675 a_14266_8900.t54 a_14266_8900.t22 113.753
R676 a_14266_8900.t54 a_14266_8900.t15 113.753
R677 a_14266_8900.t54 a_14266_8900.t33 113.753
R678 a_14266_8900.t54 a_14266_8900.t44 113.753
R679 a_14266_8900.t47 a_14266_8900.t38 113.753
R680 a_14266_8900.t47 a_14266_8900.t12 113.753
R681 a_14266_8900.t47 a_14266_8900.t4 113.753
R682 a_14266_8900.t47 a_14266_8900.t28 113.753
R683 a_14266_8900.t54 a_14266_8900.t37 113.753
R684 a_14266_8900.t54 a_14266_8900.t10 113.753
R685 a_14266_8900.t54 a_14266_8900.t3 113.753
R686 a_14266_8900.t54 a_14266_8900.t26 113.753
R687 a_14266_8900.t0 a_14266_8900.n4 57.619
R688 a_14266_8900.n4 a_14266_8900.n3 43.122
R689 a_14266_8900.n3 a_14266_8900.t1 28.571
R690 a_14266_8900.n4 a_14266_8900.t16 10.022
R691 a_14266_8900.t54 a_14266_8900.n0 5.834
R692 a_14266_8900.t47 a_14266_8900.n1 2.869
R693 a_14266_8900.t54 a_14266_8900.t47 2.813
R694 a_14266_8900.t47 a_14266_8900.n2 2.586
R695 a_52052_20860.t18 a_52052_20860.n16 2527.24
R696 a_52052_20860.n8 a_52052_20860.t7 212.622
R697 a_52052_20860.n5 a_52052_20860.t16 212.622
R698 a_52052_20860.n12 a_52052_20860.n10 208.271
R699 a_52052_20860.n2 a_52052_20860.n0 208.271
R700 a_52052_20860.n14 a_52052_20860.n12 208.271
R701 a_52052_20860.n9 a_52052_20860.n8 208.271
R702 a_52052_20860.n4 a_52052_20860.n2 208.271
R703 a_52052_20860.n6 a_52052_20860.n5 208.271
R704 a_52052_20860.n7 a_52052_20860.n6 122.265
R705 a_52052_20860.n15 a_52052_20860.n14 121.297
R706 a_52052_20860.n7 a_52052_20860.n4 63.478
R707 a_52052_20860.n15 a_52052_20860.n9 63.217
R708 a_52052_20860.n16 a_52052_20860.n7 38.746
R709 a_52052_20860.n16 a_52052_20860.n15 15.694
R710 a_52052_20860.n8 a_52052_20860.t4 4.351
R711 a_52052_20860.n9 a_52052_20860.t1 4.351
R712 a_52052_20860.n5 a_52052_20860.t13 4.351
R713 a_52052_20860.n6 a_52052_20860.t10 4.351
R714 a_52052_20860.n10 a_52052_20860.t3 4.35
R715 a_52052_20860.n10 a_52052_20860.t8 4.35
R716 a_52052_20860.n11 a_52052_20860.t0 4.35
R717 a_52052_20860.n11 a_52052_20860.t6 4.35
R718 a_52052_20860.n13 a_52052_20860.t5 4.35
R719 a_52052_20860.n13 a_52052_20860.t2 4.35
R720 a_52052_20860.n0 a_52052_20860.t12 4.35
R721 a_52052_20860.n0 a_52052_20860.t17 4.35
R722 a_52052_20860.n1 a_52052_20860.t9 4.35
R723 a_52052_20860.n1 a_52052_20860.t15 4.35
R724 a_52052_20860.n3 a_52052_20860.t14 4.35
R725 a_52052_20860.n3 a_52052_20860.t11 4.35
R726 a_52052_20860.n14 a_52052_20860.n13 0.001
R727 a_52052_20860.n12 a_52052_20860.n11 0.001
R728 a_52052_20860.n4 a_52052_20860.n3 0.001
R729 a_52052_20860.n2 a_52052_20860.n1 0.001
R730 a_56334_20860.n0 a_56334_20860.t2 171.564
R731 a_56334_20860.n0 a_56334_20860.t1 171.563
R732 a_56334_20860.t0 a_56334_20860.n0 171.52
R733 a_23156_5032.n0 a_23156_5032.t0 365.308
R734 a_23156_5032.n2 a_23156_5032.t3 93.107
R735 a_23156_5032.n5 a_23156_5032.n4 75.71
R736 a_23156_5032.n3 a_23156_5032.n2 75.707
R737 a_23156_5032.n4 a_23156_5032.n3 75.707
R738 a_23156_5032.n1 a_23156_5032.n0 75.707
R739 a_23156_5032.n5 a_23156_5032.n1 75.706
R740 a_23156_5032.t6 a_23156_5032.n5 17.401
R741 a_23156_5032.n0 a_23156_5032.t4 17.401
R742 a_23156_5032.n1 a_23156_5032.t1 17.401
R743 a_23156_5032.n4 a_23156_5032.t2 17.401
R744 a_23156_5032.n3 a_23156_5032.t7 17.401
R745 a_23156_5032.n2 a_23156_5032.t5 17.401
R746 vbiasr.n17 vbiasr.t20 11.266
R747 vbiasr.n28 vbiasr.t32 7.425
R748 vbiasr.n17 vbiasr.t37 7.425
R749 vbiasr.n26 vbiasr.t28 5.713
R750 vbiasr.n26 vbiasr.t36 5.713
R751 vbiasr.n9 vbiasr.t35 5.713
R752 vbiasr.n9 vbiasr.t23 5.713
R753 vbiasr.n10 vbiasr.t27 5.713
R754 vbiasr.n10 vbiasr.t25 5.713
R755 vbiasr.n11 vbiasr.t34 5.713
R756 vbiasr.n11 vbiasr.t33 5.713
R757 vbiasr.n12 vbiasr.t21 5.713
R758 vbiasr.n12 vbiasr.t40 5.713
R759 vbiasr.n13 vbiasr.t24 5.713
R760 vbiasr.n13 vbiasr.t31 5.713
R761 vbiasr.n15 vbiasr.t38 5.713
R762 vbiasr.n15 vbiasr.t22 5.713
R763 vbiasr.n16 vbiasr.t29 5.713
R764 vbiasr.n16 vbiasr.t26 5.713
R765 vbiasr.n14 vbiasr.t30 5.713
R766 vbiasr.n14 vbiasr.t39 5.713
R767 vbiasr.n39 vbiasr.t12 5.244
R768 vbiasr.n29 vbiasr.t0 5.244
R769 vbiasr.n0 vbiasr.t18 3.48
R770 vbiasr.n0 vbiasr.t16 3.48
R771 vbiasr.n1 vbiasr.t3 3.48
R772 vbiasr.n1 vbiasr.t5 3.48
R773 vbiasr.n2 vbiasr.t10 3.48
R774 vbiasr.n2 vbiasr.t15 3.48
R775 vbiasr.n3 vbiasr.t14 3.48
R776 vbiasr.n3 vbiasr.t1 3.48
R777 vbiasr.n4 vbiasr.t4 3.48
R778 vbiasr.n4 vbiasr.t9 3.48
R779 vbiasr.n5 vbiasr.t8 3.48
R780 vbiasr.n5 vbiasr.t13 3.48
R781 vbiasr.n6 vbiasr.t19 3.48
R782 vbiasr.n6 vbiasr.t2 3.48
R783 vbiasr.n7 vbiasr.t7 3.48
R784 vbiasr.n7 vbiasr.t6 3.48
R785 vbiasr.n8 vbiasr.t11 3.48
R786 vbiasr.n8 vbiasr.t17 3.48
R787 vbiasr.n35 vbiasr.n3 1.766
R788 vbiasr.n38 vbiasr.n0 1.766
R789 vbiasr.n32 vbiasr.n6 1.766
R790 vbiasr.n31 vbiasr.n7 1.764
R791 vbiasr.n34 vbiasr.n4 1.762
R792 vbiasr.n36 vbiasr.n2 1.761
R793 vbiasr.n33 vbiasr.n5 1.758
R794 vbiasr.n37 vbiasr.n1 1.758
R795 vbiasr.n30 vbiasr.n8 1.754
R796 vbiasr.n21 vbiasr.n13 1.714
R797 vbiasr.n18 vbiasr.n16 1.714
R798 vbiasr.n24 vbiasr.n10 1.714
R799 vbiasr.n25 vbiasr.n9 1.712
R800 vbiasr.n22 vbiasr.n12 1.71
R801 vbiasr.n20 vbiasr.n14 1.709
R802 vbiasr.n23 vbiasr.n11 1.706
R803 vbiasr.n19 vbiasr.n15 1.706
R804 vbiasr.n27 vbiasr.n26 1.702
R805 vbiasr.n29 vbiasr.n28 0.293
R806 vbiasr vbiasr.n39 0.273
R807 vbiasr.n23 vbiasr.n22 0.031
R808 vbiasr.n34 vbiasr.n33 0.031
R809 vbiasr.n37 vbiasr.n36 0.031
R810 vbiasr.n20 vbiasr.n19 0.031
R811 vbiasr.n31 vbiasr.n30 0.031
R812 vbiasr.n27 vbiasr.n25 0.031
R813 vbiasr.n28 vbiasr.n27 0.031
R814 vbiasr.n30 vbiasr.n29 0.031
R815 vbiasr.n38 vbiasr.n37 0.03
R816 vbiasr.n19 vbiasr.n18 0.03
R817 vbiasr.n18 vbiasr.n17 0.03
R818 vbiasr.n39 vbiasr.n38 0.03
R819 vbiasr.n25 vbiasr.n24 0.03
R820 vbiasr.n32 vbiasr.n31 0.03
R821 vbiasr.n35 vbiasr.n34 0.03
R822 vbiasr.n22 vbiasr.n21 0.03
R823 vbiasr.n36 vbiasr.n35 0.03
R824 vbiasr.n21 vbiasr.n20 0.03
R825 vbiasr.n33 vbiasr.n32 0.03
R826 vbiasr.n24 vbiasr.n23 0.03
R827 a_23436_16644.t46 a_23436_16644.t43 1273.78
R828 a_23436_16644.n3 a_23436_16644.t1 1158.7
R829 a_23436_16644.n3 a_23436_16644.t60 169.095
R830 a_23436_16644.t60 a_23436_16644.t45 113.753
R831 a_23436_16644.t60 a_23436_16644.t5 113.753
R832 a_23436_16644.t60 a_23436_16644.t21 113.753
R833 a_23436_16644.t60 a_23436_16644.t20 113.753
R834 a_23436_16644.t60 a_23436_16644.t2 113.753
R835 a_23436_16644.t60 a_23436_16644.t17 113.753
R836 a_23436_16644.t60 a_23436_16644.t37 113.753
R837 a_23436_16644.t60 a_23436_16644.t33 113.753
R838 a_23436_16644.n2 a_23436_16644.t44 113.753
R839 a_23436_16644.n2 a_23436_16644.t59 113.753
R840 a_23436_16644.n2 a_23436_16644.t14 113.753
R841 a_23436_16644.n2 a_23436_16644.t32 113.753
R842 a_23436_16644.n0 a_23436_16644.t10 113.753
R843 a_23436_16644.n0 a_23436_16644.t28 113.753
R844 a_23436_16644.n1 a_23436_16644.t26 113.753
R845 a_23436_16644.n1 a_23436_16644.t34 113.753
R846 a_23436_16644.n1 a_23436_16644.t47 113.753
R847 a_23436_16644.n1 a_23436_16644.t6 113.753
R848 a_23436_16644.n1 a_23436_16644.t24 113.753
R849 a_23436_16644.n0 a_23436_16644.t50 113.753
R850 a_23436_16644.n0 a_23436_16644.t22 113.753
R851 a_23436_16644.n0 a_23436_16644.t40 113.753
R852 a_23436_16644.n0 a_23436_16644.t58 113.753
R853 a_23436_16644.t12 a_23436_16644.t56 113.753
R854 a_23436_16644.t12 a_23436_16644.t8 113.753
R855 a_23436_16644.t12 a_23436_16644.t18 113.753
R856 a_23436_16644.t12 a_23436_16644.t38 113.753
R857 a_23436_16644.t12 a_23436_16644.t54 113.753
R858 a_23436_16644.n0 a_23436_16644.t11 113.753
R859 a_23436_16644.t12 a_23436_16644.t29 113.753
R860 a_23436_16644.t12 a_23436_16644.t27 113.753
R861 a_23436_16644.t12 a_23436_16644.t35 113.753
R862 a_23436_16644.t12 a_23436_16644.t48 113.753
R863 a_23436_16644.t12 a_23436_16644.t7 113.753
R864 a_23436_16644.t12 a_23436_16644.t25 113.753
R865 a_23436_16644.n0 a_23436_16644.t51 113.753
R866 a_23436_16644.n0 a_23436_16644.t23 113.753
R867 a_23436_16644.n0 a_23436_16644.t41 113.753
R868 a_23436_16644.t12 a_23436_16644.t61 113.753
R869 a_23436_16644.t12 a_23436_16644.t57 113.753
R870 a_23436_16644.t12 a_23436_16644.t9 113.753
R871 a_23436_16644.t12 a_23436_16644.t19 113.753
R872 a_23436_16644.t12 a_23436_16644.t39 113.753
R873 a_23436_16644.t12 a_23436_16644.t55 113.753
R874 a_23436_16644.t60 a_23436_16644.t15 113.753
R875 a_23436_16644.t60 a_23436_16644.t36 113.753
R876 a_23436_16644.t60 a_23436_16644.t53 113.753
R877 a_23436_16644.t60 a_23436_16644.t52 113.753
R878 a_23436_16644.t12 a_23436_16644.t4 113.753
R879 a_23436_16644.t12 a_23436_16644.t13 113.753
R880 a_23436_16644.t12 a_23436_16644.t31 113.753
R881 a_23436_16644.t12 a_23436_16644.t49 113.753
R882 a_23436_16644.t60 a_23436_16644.t30 113.753
R883 a_23436_16644.t60 a_23436_16644.t42 113.753
R884 a_23436_16644.t60 a_23436_16644.t3 113.753
R885 a_23436_16644.t60 a_23436_16644.t16 113.753
R886 a_23436_16644.t0 a_23436_16644.n3 59.624
R887 a_23436_16644.t60 a_23436_16644.t46 6.578
R888 a_23436_16644.t60 a_23436_16644.n0 5.834
R889 a_23436_16644.t12 a_23436_16644.n1 2.869
R890 a_23436_16644.t12 a_23436_16644.n2 2.586
R891 a_23436_16644.t60 a_23436_16644.t12 2.576
R892 a_25778_4988.n0 a_25778_4988.t7 334.707
R893 a_25778_4988.n4 a_25778_4988.t2 93.107
R894 a_25778_4988.n5 a_25778_4988.n4 75.71
R895 a_25778_4988.n3 a_25778_4988.n2 75.707
R896 a_25778_4988.n2 a_25778_4988.n1 75.707
R897 a_25778_4988.n1 a_25778_4988.n0 75.707
R898 a_25778_4988.n5 a_25778_4988.n3 75.706
R899 a_25778_4988.t6 a_25778_4988.n5 17.401
R900 a_25778_4988.n0 a_25778_4988.t3 17.401
R901 a_25778_4988.n1 a_25778_4988.t0 17.401
R902 a_25778_4988.n2 a_25778_4988.t5 17.401
R903 a_25778_4988.n3 a_25778_4988.t1 17.401
R904 a_25778_4988.n4 a_25778_4988.t4 17.401
R905 Fvco.t28 Fvco.t8 1273.78
R906 Fvco.t28 Fvco.n3 132.569
R907 Fvco.t4 Fvco.t25 113.753
R908 Fvco.t4 Fvco.t24 113.753
R909 Fvco.t4 Fvco.t35 113.753
R910 Fvco.t4 Fvco.t48 113.753
R911 Fvco.n2 Fvco.t47 113.753
R912 Fvco.n2 Fvco.t23 113.753
R913 Fvco.n2 Fvco.t20 113.753
R914 Fvco.n2 Fvco.t30 113.753
R915 Fvco.n0 Fvco.t13 113.753
R916 Fvco.n0 Fvco.t27 113.753
R917 Fvco.t26 Fvco.t38 113.753
R918 Fvco.t26 Fvco.t32 113.753
R919 Fvco.t26 Fvco.t11 113.753
R920 Fvco.t26 Fvco.t6 113.753
R921 Fvco.t26 Fvco.t21 113.753
R922 Fvco.n0 Fvco.t17 113.753
R923 Fvco.n0 Fvco.t44 113.753
R924 Fvco.n0 Fvco.t42 113.753
R925 Fvco.n0 Fvco.t2 113.753
R926 Fvco.t26 Fvco.t15 113.753
R927 Fvco.t26 Fvco.t9 113.753
R928 Fvco.t26 Fvco.t40 113.753
R929 Fvco.t26 Fvco.t36 113.753
R930 Fvco.t26 Fvco.t49 113.753
R931 Fvco.n0 Fvco.t14 113.753
R932 Fvco.t26 Fvco.t29 113.753
R933 Fvco.t26 Fvco.t39 113.753
R934 Fvco.t26 Fvco.t33 113.753
R935 Fvco.t26 Fvco.t12 113.753
R936 Fvco.t26 Fvco.t7 113.753
R937 Fvco.t26 Fvco.t22 113.753
R938 Fvco.n0 Fvco.t18 113.753
R939 Fvco.n0 Fvco.t45 113.753
R940 Fvco.n0 Fvco.t43 113.753
R941 Fvco.n1 Fvco.t3 113.753
R942 Fvco.n1 Fvco.t16 113.753
R943 Fvco.n1 Fvco.t10 113.753
R944 Fvco.n1 Fvco.t41 113.753
R945 Fvco.t26 Fvco.t37 113.753
R946 Fvco.t26 Fvco.t50 113.753
R947 Fvco.t4 Fvco.t5 113.753
R948 Fvco.t4 Fvco.t34 113.753
R949 Fvco.t4 Fvco.t31 113.753
R950 Fvco.t4 Fvco.t46 113.753
R951 Fvco.t4 Fvco.t19 113.753
R952 Fvco.n3 Fvco.t0 77.367
R953 Fvco.n3 Fvco.t1 28.578
R954 Fvco.t28 Fvco.t4 5.352
R955 Fvco.t4 Fvco.t26 4.314
R956 Fvco.t4 Fvco.n0 3.605
R957 Fvco.t26 Fvco.n1 2.943
R958 Fvco.t4 Fvco.n2 2.578
R959 vbiasob.n2 vbiasob.t1 67.964
R960 vbiasob.n0 vbiasob.t3 61.399
R961 vbiasob.n0 vbiasob.t4 60.299
R962 vbiasob.n1 vbiasob.t0 18.573
R963 vbiasob.n3 vbiasob.n2 12.525
R964 vbiasob.n1 vbiasob.t2 5.717
R965 vbiasob.n2 vbiasob.n1 1.012
R966 vbiasob.n3 vbiasob.n0 0.614
R967 vbiasob vbiasob.n3 0.484
R968 a_56272_15934.t0 a_56272_15934.t1 409.924
R969 vbiasbuffer.n0 vbiasbuffer.t1 136.915
R970 vbiasbuffer.n1 vbiasbuffer.t4 125.304
R971 vbiasbuffer.n1 vbiasbuffer.t3 120.586
R972 vbiasbuffer.n0 vbiasbuffer.t0 22.405
R973 vbiasbuffer vbiasbuffer.n0 15.01
R974 vbiasbuffer.n0 vbiasbuffer.t2 5.719
R975 vbiasbuffer vbiasbuffer.n1 0.631
R976 a_57726_5786.n0 a_57726_5786.t2 85.561
R977 a_57726_5786.n1 a_57726_5786.t0 85.561
R978 a_57726_5786.n0 a_57726_5786.t5 39.685
R979 a_57726_5786.n1 a_57726_5786.t4 17.517
R980 a_57726_5786.t3 a_57726_5786.n3 5.8
R981 a_57726_5786.n3 a_57726_5786.t1 5.8
R982 a_57726_5786.n3 a_57726_5786.n2 0.736
R983 a_57726_5786.n2 a_57726_5786.n0 0.231
R984 a_57726_5786.n2 a_57726_5786.n1 0.206
R985 a_28578_5014.n5 a_28578_5014.t7 265.844
R986 a_28578_5014.n0 a_28578_5014.t5 93.107
R987 a_28578_5014.n5 a_28578_5014.n4 75.71
R988 a_28578_5014.n1 a_28578_5014.n0 75.707
R989 a_28578_5014.n2 a_28578_5014.n1 75.707
R990 a_28578_5014.n3 a_28578_5014.n2 75.707
R991 a_28578_5014.n4 a_28578_5014.n3 75.707
R992 a_28578_5014.t6 a_28578_5014.n5 17.401
R993 a_28578_5014.n4 a_28578_5014.t3 17.401
R994 a_28578_5014.n3 a_28578_5014.t1 17.401
R995 a_28578_5014.n2 a_28578_5014.t4 17.401
R996 a_28578_5014.n1 a_28578_5014.t2 17.401
R997 a_28578_5014.n0 a_28578_5014.t0 17.401
R998 CLK_BY_4_IPH_BAR.n0 CLK_BY_4_IPH_BAR.t7 458.51
R999 CLK_BY_4_IPH_BAR.n0 CLK_BY_4_IPH_BAR.t3 402.739
R1000 CLK_BY_4_IPH_BAR.n4 CLK_BY_4_IPH_BAR.t4 333.651
R1001 CLK_BY_4_IPH_BAR.n4 CLK_BY_4_IPH_BAR.t5 297.233
R1002 CLK_BY_4_IPH_BAR.n1 CLK_BY_4_IPH_BAR.t6 286.172
R1003 CLK_BY_4_IPH_BAR.n1 CLK_BY_4_IPH_BAR.t2 227.612
R1004 CLK_BY_4_IPH_BAR.n2 CLK_BY_4_IPH_BAR.n1 202.215
R1005 CLK_BY_4_IPH_BAR.n3 CLK_BY_4_IPH_BAR.n2 73.86
R1006 CLK_BY_4_IPH_BAR.t1 CLK_BY_4_IPH_BAR.n4 70.234
R1007 CLK_BY_4_IPH_BAR.n2 CLK_BY_4_IPH_BAR.n0 44.559
R1008 CLK_BY_4_IPH_BAR.n3 CLK_BY_4_IPH_BAR.t0 24.347
R1009 CLK_BY_4_IPH_BAR.t1 CLK_BY_4_IPH_BAR.n3 1.282
R1010 a_50583_13108.n0 a_50583_13108.t1 1776.66
R1011 a_50583_13108.n0 a_50583_13108.t2 171.607
R1012 a_50583_13108.t0 a_50583_13108.n0 171.607
R1013 a_27762_11446.t11 a_27762_11446.t48 1273.78
R1014 a_27762_11446.t47 a_27762_11446.t13 113.753
R1015 a_27762_11446.t47 a_27762_11446.t23 113.753
R1016 a_27762_11446.t47 a_27762_11446.t39 113.753
R1017 a_27762_11446.t47 a_27762_11446.t56 113.753
R1018 a_27762_11446.t47 a_27762_11446.t45 113.753
R1019 a_27762_11446.t47 a_27762_11446.t60 113.753
R1020 a_27762_11446.t47 a_27762_11446.t9 113.753
R1021 a_27762_11446.t47 a_27762_11446.t30 113.753
R1022 a_27762_11446.n2 a_27762_11446.t25 113.753
R1023 a_27762_11446.n2 a_27762_11446.t37 113.753
R1024 a_27762_11446.n2 a_27762_11446.t53 113.753
R1025 a_27762_11446.n2 a_27762_11446.t7 113.753
R1026 a_27762_11446.n0 a_27762_11446.t28 113.753
R1027 a_27762_11446.n0 a_27762_11446.t41 113.753
R1028 a_27762_11446.n1 a_27762_11446.t58 113.753
R1029 a_27762_11446.n1 a_27762_11446.t51 113.753
R1030 a_27762_11446.n1 a_27762_11446.t5 113.753
R1031 a_27762_11446.n1 a_27762_11446.t20 113.753
R1032 a_27762_11446.n1 a_27762_11446.t35 113.753
R1033 a_27762_11446.n0 a_27762_11446.t15 113.753
R1034 a_27762_11446.n0 a_27762_11446.t46 113.753
R1035 a_27762_11446.n0 a_27762_11446.t61 113.753
R1036 a_27762_11446.n0 a_27762_11446.t10 113.753
R1037 a_27762_11446.t21 a_27762_11446.t31 113.753
R1038 a_27762_11446.t21 a_27762_11446.t26 113.753
R1039 a_27762_11446.t21 a_27762_11446.t38 113.753
R1040 a_27762_11446.t21 a_27762_11446.t54 113.753
R1041 a_27762_11446.t21 a_27762_11446.t8 113.753
R1042 a_27762_11446.n0 a_27762_11446.t29 113.753
R1043 a_27762_11446.t21 a_27762_11446.t42 113.753
R1044 a_27762_11446.t21 a_27762_11446.t59 113.753
R1045 a_27762_11446.t21 a_27762_11446.t52 113.753
R1046 a_27762_11446.t21 a_27762_11446.t6 113.753
R1047 a_27762_11446.t21 a_27762_11446.t22 113.753
R1048 a_27762_11446.t21 a_27762_11446.t36 113.753
R1049 a_27762_11446.n0 a_27762_11446.t16 113.753
R1050 a_27762_11446.n0 a_27762_11446.t3 113.753
R1051 a_27762_11446.n0 a_27762_11446.t17 113.753
R1052 a_27762_11446.t21 a_27762_11446.t32 113.753
R1053 a_27762_11446.t21 a_27762_11446.t44 113.753
R1054 a_27762_11446.t21 a_27762_11446.t43 113.753
R1055 a_27762_11446.t21 a_27762_11446.t55 113.753
R1056 a_27762_11446.t21 a_27762_11446.t12 113.753
R1057 a_27762_11446.t21 a_27762_11446.t24 113.753
R1058 a_27762_11446.t47 a_27762_11446.t14 113.753
R1059 a_27762_11446.t47 a_27762_11446.t27 113.753
R1060 a_27762_11446.t47 a_27762_11446.t40 113.753
R1061 a_27762_11446.t47 a_27762_11446.t57 113.753
R1062 a_27762_11446.t21 a_27762_11446.t50 113.753
R1063 a_27762_11446.t21 a_27762_11446.t4 113.753
R1064 a_27762_11446.t21 a_27762_11446.t19 113.753
R1065 a_27762_11446.t21 a_27762_11446.t34 113.753
R1066 a_27762_11446.t47 a_27762_11446.t49 113.753
R1067 a_27762_11446.t47 a_27762_11446.t2 113.753
R1068 a_27762_11446.t47 a_27762_11446.t18 113.753
R1069 a_27762_11446.t47 a_27762_11446.t33 113.753
R1070 a_27762_11446.n4 a_27762_11446.n3 88.886
R1071 a_27762_11446.n4 a_27762_11446.t0 81.996
R1072 a_27762_11446.t1 a_27762_11446.n4 59.267
R1073 a_27762_11446.t47 a_27762_11446.n0 5.834
R1074 a_27762_11446.n3 a_27762_11446.t11 4.994
R1075 a_27762_11446.n3 a_27762_11446.t47 4.809
R1076 a_27762_11446.t21 a_27762_11446.n1 2.869
R1077 a_27762_11446.t47 a_27762_11446.t21 2.8
R1078 a_27762_11446.t21 a_27762_11446.n2 2.586
R1079 a_49932_4124.t1 a_49932_4124.t2 33.597
R1080 a_49932_4124.t0 a_49932_4124.t1 13.614
R1081 a_49932_4124.t1 a_49932_4124.t3 11.692
R1082 a_44752_16348.t2 a_44752_16348.n2 349.137
R1083 a_44752_16348.n1 a_44752_16348.t1 197.553
R1084 a_44752_16348.n0 a_44752_16348.t3 178.539
R1085 a_44752_16348.n0 a_44752_16348.t4 122.603
R1086 a_44752_16348.n1 a_44752_16348.t0 114.713
R1087 a_44752_16348.n2 a_44752_16348.n0 95.215
R1088 a_44752_16348.n2 a_44752_16348.n1 26.034
R1089 a_51138_19904.t0 a_51138_19904.n0 171.568
R1090 a_51138_19904.n0 a_51138_19904.t2 171.564
R1091 a_51138_19904.n0 a_51138_19904.t1 171.52
R1092 a_14832_12082.n1 a_14832_12082.t3 434.515
R1093 a_14832_12082.n0 a_14832_12082.t2 217.163
R1094 a_14832_12082.t1 a_14832_12082.n1 52.152
R1095 a_14832_12082.n0 a_14832_12082.t0 3.106
R1096 a_14832_12082.n1 a_14832_12082.n0 0.908
R1097 a_23160_10936.n5 a_23160_10936.t7 391.966
R1098 a_23160_10936.n0 a_23160_10936.t5 93.107
R1099 a_23160_10936.n5 a_23160_10936.n4 75.709
R1100 a_23160_10936.n1 a_23160_10936.n0 75.707
R1101 a_23160_10936.n2 a_23160_10936.n1 75.707
R1102 a_23160_10936.n3 a_23160_10936.n2 75.707
R1103 a_23160_10936.n4 a_23160_10936.n3 75.707
R1104 a_23160_10936.t6 a_23160_10936.n5 17.401
R1105 a_23160_10936.n4 a_23160_10936.t2 17.401
R1106 a_23160_10936.n3 a_23160_10936.t0 17.401
R1107 a_23160_10936.n2 a_23160_10936.t3 17.401
R1108 a_23160_10936.n1 a_23160_10936.t1 17.401
R1109 a_23160_10936.n0 a_23160_10936.t4 17.401
R1110 a_28438_10874.n0 a_28438_10874.t7 338.927
R1111 a_28438_10874.n4 a_28438_10874.t3 93.107
R1112 a_28438_10874.n5 a_28438_10874.n4 75.71
R1113 a_28438_10874.n1 a_28438_10874.n0 75.708
R1114 a_28438_10874.n3 a_28438_10874.n2 75.707
R1115 a_28438_10874.n2 a_28438_10874.n1 75.707
R1116 a_28438_10874.n5 a_28438_10874.n3 75.706
R1117 a_28438_10874.t6 a_28438_10874.n5 17.401
R1118 a_28438_10874.n0 a_28438_10874.t4 17.401
R1119 a_28438_10874.n1 a_28438_10874.t0 17.401
R1120 a_28438_10874.n2 a_28438_10874.t5 17.401
R1121 a_28438_10874.n3 a_28438_10874.t1 17.401
R1122 a_28438_10874.n4 a_28438_10874.t2 17.401
R1123 a_14910_6932.n1 a_14910_6932.t3 434.494
R1124 a_14910_6932.n0 a_14910_6932.t2 217.163
R1125 a_14910_6932.t1 a_14910_6932.n1 52.318
R1126 a_14910_6932.n0 a_14910_6932.t0 3.106
R1127 a_14910_6932.n1 a_14910_6932.n0 0.906
R1128 a_26016_10878.n5 a_26016_10878.t7 305.609
R1129 a_26016_10878.n0 a_26016_10878.t5 93.107
R1130 a_26016_10878.n5 a_26016_10878.n4 75.71
R1131 a_26016_10878.n1 a_26016_10878.n0 75.707
R1132 a_26016_10878.n2 a_26016_10878.n1 75.707
R1133 a_26016_10878.n3 a_26016_10878.n2 75.707
R1134 a_26016_10878.n4 a_26016_10878.n3 75.707
R1135 a_26016_10878.t6 a_26016_10878.n5 17.401
R1136 a_26016_10878.n4 a_26016_10878.t2 17.401
R1137 a_26016_10878.n3 a_26016_10878.t0 17.401
R1138 a_26016_10878.n2 a_26016_10878.t3 17.401
R1139 a_26016_10878.n1 a_26016_10878.t1 17.401
R1140 a_26016_10878.n0 a_26016_10878.t4 17.401
R1141 CLK_BY_4_IPH.n0 CLK_BY_4_IPH.t2 447.785
R1142 CLK_BY_4_IPH.n0 CLK_BY_4_IPH.t4 402.739
R1143 CLK_BY_4_IPH.n2 CLK_BY_4_IPH.t5 227.612
R1144 CLK_BY_4_IPH.n1 CLK_BY_4_IPH.t3 227.612
R1145 CLK_BY_4_IPH.n3 CLK_BY_4_IPH.n2 219.546
R1146 CLK_BY_4_IPH.n1 CLK_BY_4_IPH.n0 184.362
R1147 CLK_BY_4_IPH.n3 CLK_BY_4_IPH.t0 91.574
R1148 CLK_BY_4_IPH.n2 CLK_BY_4_IPH.n1 51.123
R1149 CLK_BY_4_IPH.n4 CLK_BY_4_IPH.t1 40.317
R1150 CLK_BY_4_IPH CLK_BY_4_IPH.n4 11.83
R1151 CLK_BY_4_IPH.n4 CLK_BY_4_IPH.n3 0.33
R1152 a_54448_7822.t0 a_54448_7822.t1 184.89
R1153 a_24410_25128.n1 a_24410_25128.t3 434.509
R1154 a_24410_25128.n0 a_24410_25128.t2 217.163
R1155 a_24410_25128.t1 a_24410_25128.n1 52.459
R1156 a_24410_25128.n0 a_24410_25128.t0 3.106
R1157 a_24410_25128.n1 a_24410_25128.n0 0.899
R1158 a_23308_802.n1 a_23308_802.t2 434.515
R1159 a_23308_802.n0 a_23308_802.t3 217.163
R1160 a_23308_802.t1 a_23308_802.n1 52.152
R1161 a_23308_802.n0 a_23308_802.t0 3.106
R1162 a_23308_802.n1 a_23308_802.n0 0.908
R1163 a_32948_24994.n1 a_32948_24994.t3 434.487
R1164 a_32948_24994.n0 a_32948_24994.t2 217.163
R1165 a_32948_24994.t1 a_32948_24994.n1 52.153
R1166 a_32948_24994.n0 a_32948_24994.t0 3.106
R1167 a_32948_24994.n1 a_32948_24994.n0 0.887
R1168 a_28790_25040.n1 a_28790_25040.t3 434.517
R1169 a_28790_25040.n0 a_28790_25040.t2 217.163
R1170 a_28790_25040.t1 a_28790_25040.n1 52.317
R1171 a_28790_25040.n0 a_28790_25040.t0 3.106
R1172 a_28790_25040.n1 a_28790_25040.n0 0.907
R1173 z.n4 z.n3 463.355
R1174 z z.n4 20.186
R1175 z.n0 z.t4 8.766
R1176 z.n2 z.t6 8.705
R1177 z.n0 z.t7 8.7
R1178 z.n0 z.t5 8.7
R1179 z.n1 z.t3 8.7
R1180 z.n1 z.t2 8.7
R1181 z.n3 z.t1 5.713
R1182 z.n3 z.t0 5.713
R1183 z.n2 z.n0 0.137
R1184 z.n2 z.n1 0.121
R1185 z.n4 z.n2 0.093
R1186 a_51532_4150.n1 a_51532_4150.t3 19.231
R1187 a_51532_4150.n0 a_51532_4150.t1 17.234
R1188 a_51532_4150.n2 a_51532_4150.t4 14.994
R1189 a_51532_4150.n0 a_51532_4150.t0 14.151
R1190 a_51532_4150.n1 a_51532_4150.t5 13.856
R1191 a_51532_4150.t2 a_51532_4150.n0 7.827
R1192 a_51532_4150.n1 a_51532_4150.n2 5.632
R1193 a_51532_4150.n2 a_51532_4150.t6 3.653
R1194 a_51532_4150.n0 a_51532_4150.n1 3.447
R1195 a_50032_16080.t0 a_50032_16080.t1 414.247
R1196 a_50511_16072.n4 a_50511_16072.n3 524.893
R1197 a_50511_16072.n4 a_50511_16072.t8 256.935
R1198 a_50511_16072.t5 a_50511_16072.n1 8.763
R1199 a_50511_16072.n2 a_50511_16072.t0 8.705
R1200 a_50511_16072.n1 a_50511_16072.t1 8.7
R1201 a_50511_16072.n1 a_50511_16072.t2 8.7
R1202 a_50511_16072.n0 a_50511_16072.t3 8.7
R1203 a_50511_16072.n0 a_50511_16072.t4 8.7
R1204 a_50511_16072.n3 a_50511_16072.t7 5.844
R1205 a_50511_16072.n3 a_50511_16072.t6 5.744
R1206 a_50511_16072.t8 a_50511_16072.t9 1.22
R1207 a_50511_16072.n1 a_50511_16072.n0 0.137
R1208 a_50511_16072.n0 a_50511_16072.n2 0.133
R1209 a_50511_16072.n0 a_50511_16072.n4 0.122
R1210 a_38070_8852.n1 a_38070_8852.t3 434.515
R1211 a_38070_8852.n0 a_38070_8852.t2 217.163
R1212 a_38070_8852.t1 a_38070_8852.n1 52.152
R1213 a_38070_8852.n0 a_38070_8852.t0 3.106
R1214 a_38070_8852.n1 a_38070_8852.n0 0.908
R1215 a_30384_802.n1 a_30384_802.t3 434.478
R1216 a_30384_802.n0 a_30384_802.t2 217.163
R1217 a_30384_802.t1 a_30384_802.n1 52.152
R1218 a_30384_802.n0 a_30384_802.t0 3.106
R1219 a_30384_802.n1 a_30384_802.n0 0.885
R1220 a_46856_21176.t0 a_46856_21176.t1 343.213
R1221 a_51138_21494.t1 a_51138_21494.t0 501.405
R1222 a_46856_19268.n0 a_46856_19268.t0 2113.41
R1223 a_46856_19268.n0 a_46856_19268.t2 171.607
R1224 a_46856_19268.t1 a_46856_19268.n0 171.607
R1225 a_51826_16054.t0 a_51826_16054.t1 445.429
R1226 a_22972_23306.n2 a_22972_23306.t4 172.018
R1227 a_22972_23306.t0 a_22972_23306.n2 171.695
R1228 a_22972_23306.n2 a_22972_23306.n1 73.17
R1229 a_22972_23306.n1 a_22972_23306.t3 28.576
R1230 a_22972_23306.n0 a_22972_23306.t1 28.565
R1231 a_22972_23306.n0 a_22972_23306.t2 28.565
R1232 a_22972_23306.n1 a_22972_23306.n0 3.497
R1233 a_54468_7504.t0 a_54468_7504.t1 178.373
C66 vbiasr gnd 127.67fF $ **FLOATING
C67 vbiasot gnd 17.09fF
C68 a_51334_14126# gnd 5.94fF
C69 a_50320_14126# gnd 7.42fF
C70 a_56602_11692# gnd 4.81fF
C71 a_55602_11692# gnd 5.68fF
C72 a_51276_14152# gnd 3.34fF
C73 a_51636_13108# gnd 8.30fF
C74 a_51041_13108# gnd 10.28fF
C75 a_50262_14152# gnd 3.87fF
C76 vbiasob gnd 11.11fF $ **FLOATING
C77 z gnd 18.94fF $ **FLOATING
C78 a_47760_15642# gnd 2.83fF
C79 vbiasbuffer gnd 15.97fF $ **FLOATING
C80 a_43010_16058# gnd 4.05fF
C81 a_42782_16060# gnd 4.44fF
C82 a_42574_15624# gnd 5.31fF
C83 a_42550_16062# gnd 4.20fF
C84 bb gnd 13.52fF
C85 aa gnd 15.18fF
C86 b gnd 11.08fF
C87 a_77560_23350# gnd 303.47fF
C88 a gnd 8.87fF
C89 a_77242_23350# gnd 331.61fF
C90 a_77586_24654# gnd 88.66fF
C91 a_77268_24654# gnd 148.90fF
C92 Vso8b gnd 20.82fF
C93 Vso7b gnd 14.60fF
C94 a_4226_11420# gnd 8.28fF
C95 a_4288_11534# gnd 5.07fF
C96 a_4226_11612# gnd 7.54fF
C97 a_4288_11726# gnd 6.25fF
C98 a_4226_11804# gnd 7.73fF
C99 Vso5b gnd 7.67fF
C100 Vso4b gnd 47.35fF
C101 Vso6b gnd 5.87fF
C102 a_4288_11918# gnd 5.18fF
C103 a_4226_11996# gnd 8.59fF
C104 a_4288_12110# gnd 6.31fF
C105 vout gnd 5.78fF
C106 a_4226_12188# gnd 6.34fF
C107 Fvco_By4_QPH_bar gnd 26.16fF $ **FLOATING
C108 Fvco_By4_QPH gnd 37.94fF $ **FLOATING
C109 CLK_IN gnd 39.37fF
C110 Vso3b gnd 26.51fF
C111 Vso2b gnd 21.36fF
C112 Vso1b gnd 22.16fF
C113 vctrl gnd 12.38fF
C114 zz gnd 2.80fF
C115 CLK_BY_4_IPH gnd 36.30fF
C116 vinit gnd 179.15fF $ **FLOATING
C117 a_34590_30714# gnd 376.66fF
C118 a_9628_32967# gnd 376.77fF
C119 vdd gnd 5573.35fF
C120 a_54468_7504.t1 gnd 2.83fF
C121 a_22972_23306.n2 gnd 2.07fF $ **FLOATING
C122 a_46856_19268.n0 gnd 7.50fF $ **FLOATING
C123 a_51138_21494.t0 gnd 2.55fF
C124 a_51138_21494.t1 gnd 3.48fF
C125 a_30384_802.n0 gnd 3.14fF $ **FLOATING
C126 a_38070_8852.n0 gnd 3.65fF $ **FLOATING
C127 a_50511_16072.n0 gnd 2.15fF $ **FLOATING
C128 a_51532_4150.n1 gnd 3.34fF $ **FLOATING
C129 a_51532_4150.n2 gnd 3.10fF $ **FLOATING
C130 z.n0 gnd 2.27fF $ **FLOATING
C131 z.n2 gnd 2.49fF $ **FLOATING
C132 z.n4 gnd 5.27fF $ **FLOATING
C133 a_28790_25040.n0 gnd 3.75fF $ **FLOATING
C134 a_32948_24994.n0 gnd 3.11fF $ **FLOATING
C135 a_23308_802.n0 gnd 3.31fF $ **FLOATING
C136 a_24410_25128.n0 gnd 3.81fF $ **FLOATING
C137 a_54448_7822.t1 gnd 3.00fF
C138 CLK_BY_4_IPH.n3 gnd 47.47fF $ **FLOATING
C139 a_14910_6932.n0 gnd 3.12fF $ **FLOATING
C140 a_14832_12082.n0 gnd 3.86fF $ **FLOATING
C141 a_51138_19904.n0 gnd 2.56fF $ **FLOATING
C142 a_49932_4124.t1 gnd 4.56fF $ **FLOATING
C143 a_27762_11446.n0 gnd 4.61fF $ **FLOATING
C144 a_27762_11446.t47 gnd 9.32fF $ **FLOATING
C145 a_27762_11446.t21 gnd 9.31fF $ **FLOATING
C146 a_27762_11446.t11 gnd 6.97fF $ **FLOATING
C147 a_27762_11446.n3 gnd 12.17fF $ **FLOATING
C148 a_27762_11446.n4 gnd 3.93fF $ **FLOATING
C149 a_50583_13108.n0 gnd 8.05fF $ **FLOATING
C150 CLK_BY_4_IPH_BAR.n2 gnd 2.26fF $ **FLOATING
C151 CLK_BY_4_IPH_BAR.t0 gnd 4.96fF
C152 CLK_BY_4_IPH_BAR.n3 gnd 41.35fF $ **FLOATING
C153 vbiasbuffer.n0 gnd 4.69fF $ **FLOATING
C154 vbiasob.n2 gnd 5.69fF $ **FLOATING
C155 vbiasob.n3 gnd 3.40fF $ **FLOATING
C156 Fvco.n0 gnd 3.40fF $ **FLOATING
C157 Fvco.t26 gnd 5.90fF $ **FLOATING
C158 Fvco.t4 gnd 13.86fF $ **FLOATING
C159 Fvco.t28 gnd 45.10fF $ **FLOATING
C160 Fvco.n3 gnd 4.49fF $ **FLOATING
C161 a_23436_16644.n0 gnd 4.67fF $ **FLOATING
C162 a_23436_16644.t60 gnd 10.21fF $ **FLOATING
C163 a_23436_16644.t12 gnd 8.90fF $ **FLOATING
C164 a_23436_16644.t46 gnd 6.39fF $ **FLOATING
C165 a_23436_16644.n3 gnd 3.27fF $ **FLOATING
C166 vbiasr.t20 gnd 25.92fF
C167 vbiasr.n17 gnd 99.64fF $ **FLOATING
C168 vbiasr.n28 gnd 3.28fF $ **FLOATING
C169 vbiasr.n29 gnd 3.26fF $ **FLOATING
C170 vbiasr.n39 gnd 3.04fF $ **FLOATING
C171 a_56334_20860.n0 gnd 2.57fF $ **FLOATING
C172 a_52052_20860.t18 gnd 3.50fF
C173 a_14266_8900.n0 gnd 5.02fF $ **FLOATING
C174 a_14266_8900.t54 gnd 9.46fF $ **FLOATING
C175 a_14266_8900.t47 gnd 10.19fF $ **FLOATING
C176 a_14266_8900.t16 gnd 12.52fF $ **FLOATING
C177 a_14266_8900.n4 gnd 10.56fF $ **FLOATING
C178 a_17685_3840.t22 gnd 2.81fF $ **FLOATING
C179 a_17685_3840.t63 gnd 2.81fF $ **FLOATING
C180 a_17685_3840.t58 gnd 2.81fF $ **FLOATING
C181 a_17685_3840.t60 gnd 2.81fF $ **FLOATING
C182 a_17685_3840.t53 gnd 2.81fF $ **FLOATING
C183 a_17685_3840.t48 gnd 2.81fF $ **FLOATING
C184 a_17685_3840.t20 gnd 2.81fF $ **FLOATING
C185 a_17685_3840.t64 gnd 2.81fF $ **FLOATING
C186 a_17685_3840.t56 gnd 2.81fF $ **FLOATING
C187 a_17685_3840.t51 gnd 2.81fF $ **FLOATING
C188 a_17685_3840.t43 gnd 6.49fF $ **FLOATING
C189 a_17685_3840.n0 gnd 11.45fF $ **FLOATING
C190 a_17685_3840.n1 gnd 7.46fF $ **FLOATING
C191 a_17685_3840.n2 gnd 7.46fF $ **FLOATING
C192 a_17685_3840.n3 gnd 7.46fF $ **FLOATING
C193 a_17685_3840.n4 gnd 7.46fF $ **FLOATING
C194 a_17685_3840.n5 gnd 7.46fF $ **FLOATING
C195 a_17685_3840.n6 gnd 7.46fF $ **FLOATING
C196 a_17685_3840.n7 gnd 7.46fF $ **FLOATING
C197 a_17685_3840.n8 gnd 7.46fF $ **FLOATING
C198 a_17685_3840.n9 gnd 6.30fF $ **FLOATING
C199 a_17685_3840.t54 gnd 3.77fF $ **FLOATING
C200 a_17685_3840.n10 gnd 7.72fF $ **FLOATING
C201 a_17685_3840.t46 gnd 2.81fF $ **FLOATING
C202 a_17685_3840.t38 gnd 2.81fF $ **FLOATING
C203 a_17685_3840.t31 gnd 2.81fF $ **FLOATING
C204 a_17685_3840.t33 gnd 2.81fF $ **FLOATING
C205 a_17685_3840.t24 gnd 2.81fF $ **FLOATING
C206 a_17685_3840.t18 gnd 2.81fF $ **FLOATING
C207 a_17685_3840.t61 gnd 2.81fF $ **FLOATING
C208 a_17685_3840.t55 gnd 2.81fF $ **FLOATING
C209 a_17685_3840.t49 gnd 2.81fF $ **FLOATING
C210 a_17685_3840.t42 gnd 2.81fF $ **FLOATING
C211 a_17685_3840.t35 gnd 6.49fF $ **FLOATING
C212 a_17685_3840.n11 gnd 11.43fF $ **FLOATING
C213 a_17685_3840.n12 gnd 7.45fF $ **FLOATING
C214 a_17685_3840.n13 gnd 7.45fF $ **FLOATING
C215 a_17685_3840.n14 gnd 7.45fF $ **FLOATING
C216 a_17685_3840.n15 gnd 7.45fF $ **FLOATING
C217 a_17685_3840.n16 gnd 7.45fF $ **FLOATING
C218 a_17685_3840.n17 gnd 7.45fF $ **FLOATING
C219 a_17685_3840.n18 gnd 7.45fF $ **FLOATING
C220 a_17685_3840.n19 gnd 7.45fF $ **FLOATING
C221 a_17685_3840.n20 gnd 6.30fF $ **FLOATING
C222 a_17685_3840.t27 gnd 3.77fF $ **FLOATING
C223 a_17685_3840.n21 gnd 5.66fF $ **FLOATING
C224 a_17685_3840.n22 gnd 6.42fF $ **FLOATING
C225 a_17685_3840.n23 gnd 3.24fF $ **FLOATING
C226 a_17685_3840.n28 gnd 2.56fF $ **FLOATING
C227 a_17685_3840.t47 gnd 2.81fF $ **FLOATING
C228 a_17685_3840.t41 gnd 2.81fF $ **FLOATING
C229 a_17685_3840.t44 gnd 2.81fF $ **FLOATING
C230 a_17685_3840.t36 gnd 2.81fF $ **FLOATING
C231 a_17685_3840.t29 gnd 2.81fF $ **FLOATING
C232 a_17685_3840.t28 gnd 2.81fF $ **FLOATING
C233 a_17685_3840.t21 gnd 2.81fF $ **FLOATING
C234 a_17685_3840.t62 gnd 2.81fF $ **FLOATING
C235 a_17685_3840.t57 gnd 2.81fF $ **FLOATING
C236 a_17685_3840.t50 gnd 6.49fF $ **FLOATING
C237 a_17685_3840.n35 gnd 11.41fF $ **FLOATING
C238 a_17685_3840.n36 gnd 7.44fF $ **FLOATING
C239 a_17685_3840.n37 gnd 7.44fF $ **FLOATING
C240 a_17685_3840.n38 gnd 7.44fF $ **FLOATING
C241 a_17685_3840.n39 gnd 7.44fF $ **FLOATING
C242 a_17685_3840.n40 gnd 7.44fF $ **FLOATING
C243 a_17685_3840.n41 gnd 7.44fF $ **FLOATING
C244 a_17685_3840.n42 gnd 7.44fF $ **FLOATING
C245 a_17685_3840.n43 gnd 7.44fF $ **FLOATING
C246 a_17685_3840.t52 gnd 2.81fF $ **FLOATING
C247 a_17685_3840.n44 gnd 6.27fF $ **FLOATING
C248 a_17685_3840.t39 gnd 3.78fF $ **FLOATING
C249 a_17685_3840.n45 gnd 7.77fF $ **FLOATING
C250 a_17685_3840.t45 gnd 2.81fF $ **FLOATING
C251 a_17685_3840.t37 gnd 2.81fF $ **FLOATING
C252 a_17685_3840.t30 gnd 2.81fF $ **FLOATING
C253 a_17685_3840.t32 gnd 2.81fF $ **FLOATING
C254 a_17685_3840.t23 gnd 2.81fF $ **FLOATING
C255 a_17685_3840.t17 gnd 2.81fF $ **FLOATING
C256 a_17685_3840.t40 gnd 2.81fF $ **FLOATING
C257 a_17685_3840.t34 gnd 2.81fF $ **FLOATING
C258 a_17685_3840.t25 gnd 2.81fF $ **FLOATING
C259 a_17685_3840.t19 gnd 2.81fF $ **FLOATING
C260 a_17685_3840.t59 gnd 6.50fF $ **FLOATING
C261 a_17685_3840.n46 gnd 11.46fF $ **FLOATING
C262 a_17685_3840.n47 gnd 7.47fF $ **FLOATING
C263 a_17685_3840.n48 gnd 7.47fF $ **FLOATING
C264 a_17685_3840.n49 gnd 7.47fF $ **FLOATING
C265 a_17685_3840.n50 gnd 7.47fF $ **FLOATING
C266 a_17685_3840.n51 gnd 7.47fF $ **FLOATING
C267 a_17685_3840.n52 gnd 7.47fF $ **FLOATING
C268 a_17685_3840.n53 gnd 7.47fF $ **FLOATING
C269 a_17685_3840.n54 gnd 7.47fF $ **FLOATING
C270 a_17685_3840.n55 gnd 6.31fF $ **FLOATING
C271 a_17685_3840.t26 gnd 3.77fF $ **FLOATING
C272 a_17685_3840.n56 gnd 5.48fF $ **FLOATING
C273 a_17685_3840.n57 gnd 6.30fF $ **FLOATING
C274 a_17685_3840.n58 gnd 3.43fF $ **FLOATING
C275 a_17685_3840.n61 gnd 2.26fF $ **FLOATING
C276 a_25099_11445.n0 gnd 4.84fF $ **FLOATING
C277 a_25099_11445.t40 gnd 9.07fF $ **FLOATING
C278 a_25099_11445.t15 gnd 10.01fF $ **FLOATING
C279 a_25099_11445.n3 gnd 2.56fF $ **FLOATING
C280 a_25099_11445.t53 gnd 8.62fF $ **FLOATING
C281 a_25099_11445.n4 gnd 7.05fF $ **FLOATING
C282 a_26036_4988.n0 gnd 9.29fF $ **FLOATING
C283 a_26036_4988.n1 gnd 4.19fF $ **FLOATING
C284 a_26036_4988.t20 gnd 9.20fF $ **FLOATING
C285 a_26036_4988.t44 gnd 6.43fF $ **FLOATING
C286 a_26036_4988.t16 gnd 5.98fF $ **FLOATING
C287 Fvco_By4_QPH.n1 gnd 11.39fF $ **FLOATING
C288 Fvco_By4_QPH.n3 gnd 2.48fF $ **FLOATING
C289 Fvco_By4_QPH.n4 gnd 2.45fF $ **FLOATING
C290 Fvco_By4_QPH.n5 gnd 5.17fF $ **FLOATING
C291 Fvco_By4_QPH.n7 gnd 5.63fF $ **FLOATING
C292 a_49874_4150.n0 gnd 4.09fF $ **FLOATING
C293 a_49874_4150.t6 gnd 2.43fF $ **FLOATING
C294 a_49874_4150.t12 gnd 2.48fF $ **FLOATING
C295 a_49874_4150.t9 gnd 2.26fF $ **FLOATING
C296 a_14188_14050.n0 gnd 9.50fF $ **FLOATING
C297 a_14188_14050.t39 gnd 4.66fF $ **FLOATING
C298 a_14188_14050.t31 gnd 20.38fF $ **FLOATING
C299 a_14188_14050.n3 gnd 3.58fF $ **FLOATING
C300 a_14188_14050.t12 gnd 10.32fF $ **FLOATING
C301 a_14188_14050.n4 gnd 10.33fF $ **FLOATING
C302 vinit.n14 gnd 8.12fF $ **FLOATING
C303 vinit.n15 gnd 174.69fF $ **FLOATING
C304 vinit.n34 gnd 2.52fF $ **FLOATING
C305 vinit.n35 gnd 2.55fF $ **FLOATING
C306 vinit.n45 gnd 5.08fF $ **FLOATING
C307 a_26690_784.n0 gnd 3.33fF $ **FLOATING
C308 a_23414_5032.n0 gnd 7.27fF $ **FLOATING
C309 a_23414_5032.t14 gnd 13.09fF $ **FLOATING
C310 a_23414_5032.n4 gnd 2.35fF $ **FLOATING
C311 a_23414_5032.t2 gnd 6.60fF $ **FLOATING
C312 a_23414_5032.n5 gnd 5.52fF $ **FLOATING
C313 a_26368_16652.n0 gnd 4.17fF $ **FLOATING
C314 a_26368_16652.t52 gnd 11.83fF $ **FLOATING
C315 a_26368_16652.t39 gnd 8.95fF $ **FLOATING
C316 a_26368_16652.t24 gnd 5.97fF $ **FLOATING
C317 a_26368_16652.n3 gnd 4.09fF $ **FLOATING
C318 Fvco_By4_QPH_bar.n0 gnd 21.37fF $ **FLOATING
C319 Fvco_By4_QPH_bar.n2 gnd 3.86fF $ **FLOATING
C320 Fvco_By4_QPH_bar.n3 gnd 3.48fF $ **FLOATING
C321 Fvco_By4_QPH_bar.n5 gnd 7.86fF $ **FLOATING
